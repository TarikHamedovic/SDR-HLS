// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Tue Mar 19 23:07:44 2024
//
// Verilog Description of module top
//

module top (i_Rx_Serial, o_Tx_Serial, led, XOut, RFIn, DiffOut, 
            PWMOut, PWMOutP1, PWMOutP2, PWMOutP3, PWMOutP4, PWMOutN1, 
            PWMOutN2, PWMOutN3, PWMOutN4, sinGen, sin_out, CIC_out_clkSin, 
            clk_25mhz) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(45[8:11])
    input i_Rx_Serial;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(47[13:24])
    output o_Tx_Serial;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(48[11:22])
    output [7:0]led;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    output XOut;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(53[9:13])
    input RFIn;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(54[9:13])
    output DiffOut;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(55[9:16])
    output PWMOut;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(56[9:15])
    output PWMOutP1;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(57[9:17])
    output PWMOutP2;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(58[9:17])
    output PWMOutP3;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(59[9:17])
    output PWMOutP4;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(60[9:17])
    output PWMOutN1;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(61[9:17])
    output PWMOutN2;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(62[9:17])
    output PWMOutN3;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(63[9:17])
    output PWMOutN4;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(64[9:17])
    output sinGen;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(65[9:15])
    output sin_out;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(66[9:16])
    output CIC_out_clkSin;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(67[9:23])
    input clk_25mhz;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(68[8:17])
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(68[8:17])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(89[6:21])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, led_c_7, led_c_6, led_c_5, 
        led_c_4, led_c_3, led_c_2, led_c_1, led_c_0, RFIn_c, DiffOut_c, 
        PWMOutP4_c, PWMOutN4_c, sinGen_c, o_Rx_DV, o_Rx_DV1;
    wire [7:0]o_Rx_Byte1;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(80[11:21])
    wire [11:0]MixerOutSin;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(85[20:31])
    wire [11:0]MixerOutCos;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(86[20:31])
    wire [11:0]CIC1_outSin;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(88[20:31])
    wire [11:0]CIC1_outCos;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(91[20:31])
    wire [63:0]phase_accum;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(93[13:24])
    wire [12:0]LOSine;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(94[20:26])
    wire [12:0]LOCosine;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(95[20:28])
    wire [63:0]phase_inc_carrGen;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(97[19:36])
    wire [63:0]phase_inc_carrGen1;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(98[19:37])
    wire [11:0]DemodOut;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(101[20:28])
    
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire [7:0]CICGain;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(103[11:18])
    
    wire n102, n16795, n99, n96, n93, n7, n6, n5, n4, n3, 
        n2, n37, n36, n35, n34, n33, n32, n31, n30_adj_2748, 
        n29_adj_2749, n28_adj_2750, n27_adj_2751, n26_adj_2752, n25_adj_2753, 
        n24_adj_2754, n23_adj_2755, n22, n21, n20, n19, n18, n17, 
        n2586, n16794, n16, n15, n14, n13, n12, n11, n10, 
        n9, n8, n7_adj_2756, n6_adj_2757, n5_adj_2758, n4_adj_2759, 
        n3_adj_2760, n2_adj_2761, n16793, n16556, n90, n16792, n16791, 
        n2443, n16785, n16784, n16783, n16782, n16781, n16775, 
        n16774, n16773, n16772, n16771, n16770, n16764, n16763, 
        n16762, n2414, n16761, n16760, n16759, n16758, n2409, 
        n16757, n16756, n2403, n16750, n16749, n16748, n16747, 
        n16746, n16745, n16744, n16326, cout, n87, n2354;
    wire [63:0]phase_accum_adj_5665;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(29[19:30])
    
    wire n2355;
    wire [11:0]MixerOutSin_11__N_236;
    wire [11:0]MixerOutCos_11__N_250;
    wire [71:0]d_tmp;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(30[26:31])
    wire [71:0]d_d_tmp;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(30[33:40])
    wire [71:0]d1;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(35[26:28])
    wire [71:0]d2;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(36[26:28])
    wire [71:0]d3;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(37[26:28])
    wire [71:0]d4;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(38[26:28])
    wire [71:0]d5;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(39[26:28])
    wire [71:0]d6;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(43[26:28])
    wire [71:0]d_d6;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(43[30:34])
    wire [71:0]d7;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(44[26:28])
    wire [71:0]d_d7;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(44[30:34])
    wire [71:0]d8;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(45[26:28])
    wire [71:0]d_d8;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(45[30:34])
    wire [71:0]d9;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(46[26:28])
    wire [71:0]d_d9;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(46[30:34])
    
    wire n84;
    wire [15:0]count;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(50[14:19])
    wire [71:0]d1_71__N_418;
    wire [71:0]d2_71__N_490;
    wire [71:0]d3_71__N_562;
    wire [71:0]d4_71__N_634;
    wire [71:0]d5_71__N_706;
    
    wire n16743, n16336, n16742, n16741, n16740, n16739, n16738, 
        n16737, n16736, n16735, n16734, n16733, n16732, n16731, 
        n16730, n16729, n81;
    wire [71:0]d6_71__N_1459;
    wire [71:0]d7_71__N_1531;
    wire [71:0]d8_71__N_1603;
    wire [71:0]d9_71__N_1675;
    
    wire n78, n183, n180, n177, n174, n171, n168, n165, n162, 
        n159, n156, n153, n150, n147, n144, n141, n138, n135, 
        n132, n129, n126, n123, n120, n117, n114, n111, n108, 
        n105, n102_adj_2762, n99_adj_2763, n96_adj_2764, n93_adj_2765, 
        n90_adj_2766, n87_adj_2767, n84_adj_2768, n81_adj_2769, n78_adj_2770, 
        n183_adj_2771, n180_adj_2772, n177_adj_2773, n174_adj_2774, 
        n171_adj_2775, n168_adj_2776, n165_adj_2777, n162_adj_2778, 
        n159_adj_2779, n156_adj_2780, n153_adj_2781, n150_adj_2782, 
        n147_adj_2783, n144_adj_2784, n141_adj_2785, n138_adj_2786, 
        n135_adj_2787, n132_adj_2788, n129_adj_2789, n126_adj_2790, 
        n123_adj_2791, n120_adj_2792, n117_adj_2793, n114_adj_2794, 
        n111_adj_2795, n108_adj_2796, n105_adj_2797, n102_adj_2798, 
        n99_adj_2799, n96_adj_2800, n93_adj_2801, n90_adj_2802, n87_adj_2803, 
        n84_adj_2804, n81_adj_2805, n78_adj_2806, n301, n298, n295, 
        n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, 
        n238, n235, n232, n229, n226, n223, n220, n217, n214, 
        n211, n208, n205, n202, n199, n196, n193, n190, n187, 
        n184, n181, n178, n175, n172, n169, n166;
    wire [71:0]d_tmp_adj_5671;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(30[26:31])
    wire [71:0]d_d_tmp_adj_5672;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(30[33:40])
    wire [71:0]d1_adj_5673;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(35[26:28])
    wire [71:0]d2_adj_5674;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(36[26:28])
    wire [71:0]d3_adj_5675;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(37[26:28])
    wire [71:0]d4_adj_5676;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(38[26:28])
    wire [71:0]d5_adj_5677;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(39[26:28])
    wire [71:0]d6_adj_5678;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(43[26:28])
    wire [71:0]d_d6_adj_5679;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(43[30:34])
    wire [71:0]d7_adj_5680;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(44[26:28])
    wire [71:0]d_d7_adj_5681;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(44[30:34])
    wire [71:0]d8_adj_5682;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(45[26:28])
    wire [71:0]d_d8_adj_5683;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(45[30:34])
    wire [71:0]d9_adj_5684;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(46[26:28])
    wire [71:0]d_d9_adj_5685;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(46[30:34])
    wire [71:0]d10_adj_5686;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(47[26:29])
    wire [15:0]count_adj_5688;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(50[14:19])
    wire [71:0]d1_71__N_418_adj_5689;
    wire [71:0]d2_71__N_490_adj_5690;
    wire [71:0]d3_71__N_562_adj_5691;
    wire [71:0]d4_71__N_634_adj_5692;
    wire [71:0]d5_71__N_706_adj_5693;
    
    wire n16419, n16728, n16727, n16726, n16725, n16724, n16723, 
        n16722, n16721, n16720, n16719, n163, n160, n157, n154, 
        n151, n148, n145, n142, n139, n136, n133, n130, n127, 
        n124;
    wire [71:0]d6_71__N_1459_adj_5705;
    wire [71:0]d7_71__N_1531_adj_5706;
    wire [71:0]d8_71__N_1603_adj_5707;
    wire [71:0]d9_71__N_1675_adj_5708;
    
    wire n16325, n16324, n16319, n16318, n16317, n16316, n16315, 
        n16314, n16313, n16312, n16311, n16310, n16309, n16308, 
        n16307, n16306, n16305, n16304, n16303, n16302, n16298, 
        n16297, n16296, n16295, n16294, n16293;
    wire [71:0]d_out_11__N_1819_adj_5711;
    
    wire n183_adj_4551, n180_adj_4552, n177_adj_4553, n174_adj_4554, 
        n171_adj_4555, n168_adj_4556, n165_adj_4557, n162_adj_4558, 
        n159_adj_4559, n156_adj_4560, n153_adj_4561, n150_adj_4562, 
        n147_adj_4563, n16368, n321, n318, n315, n312, n309, n306, 
        n303, n300, n16552, n16551, n297, n16335, n294, n16550, 
        n291, n16549, n16548, n16547, n16546, n16545, n288, n16544, 
        n11_adj_4564, n16543, n285, n282, n279, n276, n273, n16542, 
        n270, n16541;
    wire [9:0]counter;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(7[11:18])
    wire [11:0]DataInReg;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(10[12:21])
    
    wire n267, n264, n16540, n16383;
    wire [11:0]DataInReg_11__N_1856;
    
    wire n16292, n16291;
    wire [31:0]ISquare;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(24[14:21])
    
    wire n3_adj_4565, n2_adj_4566, n16418;
    wire [23:0]MultResult1;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(30[22:33])
    wire [23:0]MultResult2;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(35[22:33])
    
    wire n21_adj_4567, n20_adj_4568, n19_adj_4569, n18_adj_4570, n17_adj_4571, 
        n16_adj_4572, n16539, n15_adj_4573, n16538, n16537, n16536, 
        n261, n16535, n10_adj_4574, n2350, n14_adj_4575, n258, n2349, 
        n2348, n13_adj_4576, n209, n2347, n2346, n255, n252, n16533, 
        n12_adj_4577, n2345, n2344, n37_adj_4578, n36_adj_4579, n35_adj_4580, 
        n34_adj_4581, n33_adj_4582, n32_adj_4583, n31_adj_4584, n30_adj_4585, 
        n29_adj_4586, n28_adj_4587, n27_adj_4588, n26_adj_4589, n249, 
        n105_adj_4590, n108_adj_4591, n11_adj_4592, n25_adj_4593, n2343, 
        n24_adj_4594, n23_adj_4595, n22_adj_4596, n21_adj_4597, n20_adj_4598, 
        n19_adj_4599, n18_adj_4600, n17_adj_4601, n16_adj_4602, n15_adj_4603, 
        n14_adj_4604, n13_adj_4605, n12_adj_4606, n11_adj_4607, n10_adj_4608, 
        n9_adj_4609, n8_adj_4610, n2342, n7_adj_4611, n6_adj_4612, 
        n5_adj_4613, n4_adj_4614, n3_adj_4615, n2_adj_4616, n16417;
    wire [17:0]d_out_d_11__N_1874;
    
    wire d_out_d_11__N_1873, n10_adj_4617, n2341, n37_adj_4618, n36_adj_4619, 
        n35_adj_4620, n34_adj_4621, n33_adj_4622, n32_adj_4623, n31_adj_4624;
    wire [17:0]d_out_d_11__N_1876;
    
    wire n246, d_out_d_11__N_1875, n9_adj_4625, n30_adj_4626, n2339, 
        n29_adj_4627, n28_adj_4628, n27_adj_4629, n26_adj_4630, n25_adj_4631, 
        n24_adj_4632, n23_adj_4633, n22_adj_4634, n21_adj_4635, n20_adj_4636, 
        n19_adj_4637, n18_adj_4638, n17_adj_4639, n16_adj_4640, n15_adj_4641, 
        n14_adj_4642, n13_adj_4643, n2338, n12_adj_4644, n11_adj_4645, 
        n10_adj_4646, n9_adj_4647, n8_adj_4648, n7_adj_4649, n6_adj_4650, 
        n5_adj_4651, n4_adj_4652, n3_adj_4653, n2_adj_4654, n16532;
    wire [17:0]d_out_d_11__N_1878;
    
    wire n243, n240, d_out_d_11__N_1877, n8_adj_4655, n2337, n2336, 
        n37_adj_4656, n36_adj_4657;
    wire [17:0]d_out_d_11__N_1880;
    
    wire n237, d_out_d_11__N_1879, n7_adj_4658, n35_adj_4659, n34_adj_4660, 
        n33_adj_4661, n32_adj_4662, n31_adj_4663, n30_adj_4664, n29_adj_4665, 
        n28_adj_4666, n27_adj_4667, n26_adj_4668, n25_adj_4669, n24_adj_4670, 
        n23_adj_4671, n22_adj_4672, n21_adj_4673, n20_adj_4674, n19_adj_4675, 
        n18_adj_4676, n2334, n17_adj_4677, n16_adj_4678, n15_adj_4679, 
        n14_adj_4680, n13_adj_4681, n9_adj_4682, n10_adj_4683, n11_adj_4684, 
        n12_adj_4685, n8_adj_4686, n234;
    wire [17:0]d_out_d_11__N_1882;
    
    wire n231, n6_adj_4687, n2333, n228, n37_adj_4688, n5_adj_4689, 
        n4_adj_4690, n3_adj_4691, n2_adj_4692, n36_adj_4693, n2332, 
        n35_adj_4694, n34_adj_4695, n33_adj_4696;
    wire [17:0]d_out_d_11__N_1884;
    
    wire n225, n16381, n16379, n16371, n16372, n16374, n16375, 
        n3720, n16377, n16346, n3716, n3715, n16384, n16385, n16387, 
        n16380, n16391, n16376, n16389, n16353, n16334, n16333, 
        n16332;
    wire [17:0]d_out_d_11__N_1886;
    
    wire n222, n16290, n16331, n16330, n16329, n16340, n16341, 
        n3685, n16347, n16378, n16348, n16349, n16531, n16350, 
        n16352, n3677, n16388, n16354, n16355, n16356, n16357, 
        n16358, n16359, n16360, n16361, n16362, n16363;
    wire [17:0]d_out_d_11__N_1888;
    
    wire n219, n16530, n37_adj_4697, n36_adj_4698, n35_adj_4699;
    wire [17:0]d_out_d_11__N_1890;
    
    wire n216, n34_adj_4700, n33_adj_4701, n32_adj_4702, n31_adj_4703, 
        n30_adj_4704, n29_adj_4705, n28_adj_4706, n27_adj_4707, n26_adj_4708, 
        n25_adj_4709, n24_adj_4710, n23_adj_4711, n22_adj_4712, n21_adj_4713, 
        n20_adj_4714, n19_adj_4715, n18_adj_4716, n17_adj_4717, n16_adj_4718, 
        n15_adj_4719, n14_adj_4720, n13_adj_4721, n12_adj_4722, n11_adj_4723, 
        n10_adj_4724, n9_adj_4725, n8_adj_4726, n7_adj_4727, n6_adj_4728, 
        n5_adj_4729, n16416;
    wire [17:0]d_out_d_11__N_1892;
    
    wire n912, n913, n914, n915, n916, n917, n918, n919, n920, 
        n921, n922, n923, n924, n925, n926, n927, n4_adj_4730;
    wire [17:0]d_out_d_11__N_2353;
    wire [17:0]d_out_d_11__N_2335;
    
    wire n2353, n16529, n16528, n16527, n16526, n2356, n16525, 
        n16524, n16523, n16289, n16_adj_4731, n213, n210, n207, 
        n2358, n16700, n16699, n16698, n16697, n16696, n16695, 
        n16694, n16693, n16692, n16288, n16522, n16521, n16520, 
        n16519, n16518, n16517, n18137, n2357, n16691, n16690, 
        n16689, n16688, n16687, n16686, n16685, n16684, n16683, 
        n16287, n16285, n16284, n16516, n16512, n16681, n16680, 
        n16679, n16678, n16677, n16676, n16283, n16282, n16281, 
        n16280, n16279, n16278, n16277, n16276, n16275, n16274, 
        n16273, n16272, n16271, n16270, n16269, n16268, n16267, 
        n16266, n16265, n204, n16511, n201, n18136, n18135, n18134, 
        n198, n195, n18150, n18149, n192, n16510, n189, n17_adj_4732, 
        n186, n16509, n16675, n16328, n183_adj_4733, n2391, n2390, 
        n2389, n2388, n2387, n2386, n2385, n2384, n2383, n2382, 
        n2380, n2379, n2378, n2377, n2376, n2375, n2374, n2372, 
        n16674, n16673, n2579, n16672, n12221, n2575, n12219, 
        n16671, n12217, n16670, n16327, n12215, n2563, n12213, 
        n16669, n16338, n16668, n12211, n16667, n2542, n12209, 
        n16666, n12207, n16665, n2536, n16664, n180_adj_4734, n177_adj_4735, 
        cout_adj_4736, n16508, n16507, n16506, n16505, n16504, n16503, 
        n16502, n16501, n16500, n16499, n16498, n16497, n16496, 
        n16495, n16494, n18191, n17963, n16662, n16493, n16661, 
        n16660, n174_adj_4737, n171_adj_4738, n144_adj_4739, n141_adj_4740, 
        n138_adj_4741, n111_adj_4742, n168_adj_4743, n114_adj_4744, 
        n117_adj_4745, n120_adj_4746, n123_adj_4747, n165_adj_4748, 
        n63, n64, n65, n66, n162_adj_4749, n18267, n159_adj_4750, 
        n156_adj_4751, n153_adj_4752, n16412, n16492, n18190, n16659, 
        n150_adj_4753, n2369, n2368, n2367, n2366, n2365, n2364, 
        n2363, n2362, n2361, n2360, n2359, n147_adj_4754, n16658, 
        n16657, n16656, n15_adj_4755, n14_adj_4756, n13_adj_4757, 
        n12_adj_4758, n11_adj_4759, n10_adj_4760, n9_adj_4761, n8_adj_4762, 
        n7_adj_4763, n6_adj_4764, n5_adj_4765, n4_adj_4766, n3_adj_4767, 
        n2_adj_4768, n16491, n144_adj_4769, n16655, n16654, n16653, 
        n16652, n16651, n16650, n16649, n16648, n16647, n2593, 
        n16564, n16646, n18189, n2451, n16645, n37_adj_4770, n36_adj_4771, 
        n35_adj_4772, n34_adj_4773, n16644, n33_adj_4774, n32_adj_4775, 
        n31_adj_4776, n30_adj_4777, n29_adj_4778, n28_adj_4779, n27_adj_4780, 
        n26_adj_4781, n25_adj_4782, n24_adj_4783, n16490, n16489, 
        n16643, n141_adj_4784, n138_adj_4785, n135_adj_4786, n132_adj_4787, 
        n126_adj_4788, n129_adj_4789, n132_adj_4790, n135_adj_4791, 
        n2845, n16642, n2446, n16264, n16263, n16488, n17319, 
        n17322, n16487, n32_adj_4792, n34_adj_4793, n33_adj_4794, 
        n32_adj_4795, n31_adj_4796, n30_adj_4797, n29_adj_4798, n28_adj_4799, 
        n27_adj_4800, n26_adj_4801, n25_adj_4802, n24_adj_4803, n23_adj_4804, 
        n22_adj_4805, n21_adj_4806, n20_adj_4807, n19_adj_4808, n18_adj_4809, 
        n35_adj_4810, n36_adj_4811, n16486, n37_adj_4812, n16485, 
        n31_adj_4813, n23_adj_4814, n22_adj_4815, n21_adj_4816, n20_adj_4817, 
        n19_adj_4818, n18_adj_4819, n17_adj_4820, n16_adj_4821, n15_adj_4822, 
        n14_adj_4823, n13_adj_4824, n12_adj_4825, n11_adj_4826, n10_adj_4827, 
        n9_adj_4828, n8_adj_4829, n7_adj_4830, n6_adj_4831, n5_adj_4832, 
        n4_adj_4833, n3_adj_4834, n2_adj_4835, n22_adj_4836, n16641, 
        n78_adj_4837, n81_adj_4838, n84_adj_4839, n87_adj_4840, n90_adj_4841, 
        n93_adj_4842, n96_adj_4843, n99_adj_4844, n102_adj_4845, n105_adj_4846, 
        n108_adj_4847, n111_adj_4848, n114_adj_4849, n117_adj_4850, 
        n120_adj_4851, n123_adj_4852, n126_adj_4853, n129_adj_4854, 
        n132_adj_4855, n135_adj_4856, n138_adj_4857, n141_adj_4858, 
        n144_adj_4859, n147_adj_4860, n150_adj_4861, n153_adj_4862, 
        n156_adj_4863, n159_adj_4864, n162_adj_4865, n165_adj_4866, 
        n168_adj_4867, n171_adj_4868, n174_adj_4869, n177_adj_4870, 
        n180_adj_4871, n183_adj_4872, n78_adj_4873, n81_adj_4874, n84_adj_4875, 
        n87_adj_4876, n90_adj_4877, n93_adj_4878, n96_adj_4879, n99_adj_4880, 
        n102_adj_4881, n105_adj_4882, n108_adj_4883, n111_adj_4884, 
        n114_adj_4885, n117_adj_4886, n120_adj_4887, n123_adj_4888, 
        n126_adj_4889, n129_adj_4890, n132_adj_4891, n135_adj_4892, 
        n138_adj_4893, n141_adj_4894, n144_adj_4895, n147_adj_4896, 
        n150_adj_4897, n153_adj_4898, n156_adj_4899, n159_adj_4900, 
        n162_adj_4901, n165_adj_4902, n168_adj_4903, n171_adj_4904, 
        n174_adj_4905, n177_adj_4906, n180_adj_4907, n183_adj_4908, 
        n78_adj_4909, n81_adj_4910, n84_adj_4911, n87_adj_4912, n90_adj_4913, 
        n93_adj_4914, n96_adj_4915, n99_adj_4916, n102_adj_4917, n105_adj_4918, 
        n108_adj_4919, n111_adj_4920, n114_adj_4921, n117_adj_4922, 
        n120_adj_4923, n78_adj_4924, n81_adj_4925, n84_adj_4926, n87_adj_4927, 
        n90_adj_4928, n93_adj_4929, n96_adj_4930, n99_adj_4931, n102_adj_4932, 
        n105_adj_4933, n108_adj_4934, n111_adj_4935, n114_adj_4936, 
        n117_adj_4937, n120_adj_4938, n123_adj_4939, n126_adj_4940, 
        n129_adj_4941, n132_adj_4942, n135_adj_4943, n138_adj_4944, 
        n141_adj_4945, n144_adj_4946, n147_adj_4947, n150_adj_4948, 
        n153_adj_4949, n156_adj_4950, n159_adj_4951, n162_adj_4952, 
        n165_adj_4953, n168_adj_4954, n171_adj_4955, n174_adj_4956, 
        n177_adj_4957, n180_adj_4958, n183_adj_4959, n78_adj_4960, n81_adj_4961, 
        n84_adj_4962, n87_adj_4963, n90_adj_4964, n93_adj_4965, n96_adj_4966, 
        n99_adj_4967, n102_adj_4968, n105_adj_4969, n108_adj_4970, n111_adj_4971, 
        n114_adj_4972, n117_adj_4973, n120_adj_4974, n123_adj_4975, 
        n126_adj_4976, n129_adj_4977, n132_adj_4978, n135_adj_4979, 
        n138_adj_4980, n141_adj_4981, n144_adj_4982, n147_adj_4983, 
        n150_adj_4984, n153_adj_4985, n156_adj_4986, n159_adj_4987, 
        n162_adj_4988, n165_adj_4989, n168_adj_4990, n171_adj_4991, 
        n174_adj_4992, n177_adj_4993, n180_adj_4994, n183_adj_4995, 
        n134, n137, n140, n143, n146, n149, n152, n155, n158, 
        n161, n164, n167, n170, n173, n176, n179, n182, n185, 
        n188, n191, n194, n197, n200, n203, n206, n209_adj_4996, 
        n212, n215, n218, n221, n224, n227, n230, n233, n236, 
        n239, n242, n245, n248, n251, n254, n257, n260, n263, 
        n266, n269, n272, n275, n278, n281, n284, n287, n290, 
        n293, n296, n299, n302, n305, n308, n311, n314, n317, 
        n320, n323, n16262, n16261, n16260, n16259, n16258, n16257, 
        n16256, n16255, n16254, n16253, cout_adj_4997, cout_adj_4998, 
        n40, n49, n78_adj_4999, n81_adj_5000, n84_adj_5001, n87_adj_5002, 
        n90_adj_5003, n93_adj_5004, n96_adj_5005, n99_adj_5006, n102_adj_5007, 
        n105_adj_5008, n108_adj_5009, n111_adj_5010, n114_adj_5011, 
        n117_adj_5012, n120_adj_5013, n123_adj_5014, n126_adj_5015, 
        n129_adj_5016, n132_adj_5017, n135_adj_5018, n138_adj_5019, 
        n141_adj_5020, n144_adj_5021, n147_adj_5022, n150_adj_5023, 
        n153_adj_5024, n156_adj_5025, n159_adj_5026, n162_adj_5027, 
        n165_adj_5028, n168_adj_5029, n171_adj_5030, n174_adj_5031, 
        n177_adj_5032, n180_adj_5033, n183_adj_5034, n78_adj_5035, n81_adj_5036, 
        n84_adj_5037, n87_adj_5038, n90_adj_5039, n93_adj_5040, n96_adj_5041, 
        n99_adj_5042, n102_adj_5043, n105_adj_5044, n108_adj_5045, n111_adj_5046, 
        n114_adj_5047, n117_adj_5048, n120_adj_5049, cout_adj_5050, 
        n78_adj_5051, n81_adj_5052, n84_adj_5053, n87_adj_5054, n90_adj_5055, 
        n93_adj_5056, n96_adj_5057, n99_adj_5058, n102_adj_5059, n105_adj_5060, 
        n108_adj_5061, n111_adj_5062, n114_adj_5063, n117_adj_5064, 
        n120_adj_5065, n123_adj_5066, n126_adj_5067, n129_adj_5068, 
        n132_adj_5069, n135_adj_5070, n138_adj_5071, n141_adj_5072, 
        n144_adj_5073, n147_adj_5074, n150_adj_5075, n153_adj_5076, 
        n156_adj_5077, n159_adj_5078, n162_adj_5079, n165_adj_5080, 
        n168_adj_5081, n171_adj_5082, n174_adj_5083, n177_adj_5084, 
        n180_adj_5085, n183_adj_5086, cout_adj_5087, cout_adj_5088, 
        cout_adj_5089, n36_adj_5090, n39, n42, n45, n48, n51, 
        n54, n57, n60, n63_adj_5091, n66_adj_5092, n69, n72, n75, 
        n78_adj_5093, n81_adj_5094, n78_adj_5095, n81_adj_5096, n84_adj_5097, 
        n87_adj_5098, n90_adj_5099, n93_adj_5100, n96_adj_5101, n99_adj_5102, 
        n102_adj_5103, n105_adj_5104, n108_adj_5105, n111_adj_5106, 
        n114_adj_5107, n117_adj_5108, n120_adj_5109, n123_adj_5110, 
        n126_adj_5111, n129_adj_5112, n132_adj_5113, n135_adj_5114, 
        n138_adj_5115, n141_adj_5116, n144_adj_5117, n147_adj_5118, 
        n150_adj_5119, n153_adj_5120, n156_adj_5121, n159_adj_5122, 
        n162_adj_5123, n165_adj_5124, n168_adj_5125, n171_adj_5126, 
        n174_adj_5127, n177_adj_5128, n180_adj_5129, n183_adj_5130, 
        cout_adj_5131, cout_adj_5132, n45_adj_5133, n48_adj_5134, n51_adj_5135, 
        n54_adj_5136, n57_adj_5137, n60_adj_5138, n63_adj_5139, n66_adj_5140, 
        n69_adj_5141, n72_adj_5142, n75_adj_5143, n78_adj_5144, n81_adj_5145, 
        n84_adj_5146, n87_adj_5147, n90_adj_5148, cout_adj_5149, cout_adj_5150, 
        n76, n79, n82, n85, n88, n91, n94, n97, n100, n103, 
        n106, n109, n112, n115, n118, n36_adj_5151, n39_adj_5152, 
        n42_adj_5153, n45_adj_5154, n48_adj_5155, n51_adj_5156, n54_adj_5157, 
        n57_adj_5158, n60_adj_5159, n63_adj_5160, n66_adj_5161, n69_adj_5162, 
        n72_adj_5163, n75_adj_5164, n78_adj_5165, n81_adj_5166, n54_adj_5167, 
        n57_adj_5168, n60_adj_5169, n63_adj_5170, n66_adj_5171, n69_adj_5172, 
        n72_adj_5173, n75_adj_5174, n78_adj_5175, n81_adj_5176, n84_adj_5177, 
        n87_adj_5178, n90_adj_5179, n93_adj_5180, n96_adj_5181, n99_adj_5182, 
        n102_adj_5183, n105_adj_5184, n108_adj_5185, n111_adj_5186, 
        n114_adj_5187, n117_adj_5188, n120_adj_5189, n123_adj_5190, 
        n126_adj_5191, cout_adj_5192, n78_adj_5193, n81_adj_5194, n84_adj_5195, 
        n87_adj_5196, n90_adj_5197, n93_adj_5198, n96_adj_5199, n99_adj_5200, 
        n102_adj_5201, n105_adj_5202, n108_adj_5203, n111_adj_5204, 
        n114_adj_5205, n117_adj_5206, n120_adj_5207, n123_adj_5208, 
        n126_adj_5209, n129_adj_5210, n132_adj_5211, n135_adj_5212, 
        n138_adj_5213, n141_adj_5214, n144_adj_5215, n147_adj_5216, 
        n150_adj_5217, n153_adj_5218, n156_adj_5219, n159_adj_5220, 
        n162_adj_5221, n165_adj_5222, n168_adj_5223, n171_adj_5224, 
        n174_adj_5225, n177_adj_5226, n180_adj_5227, n183_adj_5228, 
        n16252, n16251, n16250, n16249, n16248, n16247, n16246, 
        n16245, n16244, n16243, n16242, n16241, n16240, n16239, 
        n16238, n16237, n16236, n16235, n16234, n16233, n16232, 
        n16231, n16230, n16229, n16228, n16227, n16226, n16225, 
        n16224, n16223, n16222, n16221, n16220, n16219, n16218, 
        n16217, cout_adj_5229, cout_adj_5230, n78_adj_5231, n81_adj_5232, 
        n84_adj_5233, n87_adj_5234, n90_adj_5235, n93_adj_5236, n96_adj_5237, 
        n99_adj_5238, n102_adj_5239, n105_adj_5240, n108_adj_5241, n111_adj_5242, 
        n114_adj_5243, n117_adj_5244, n120_adj_5245, n123_adj_5246, 
        n126_adj_5247, n129_adj_5248, n132_adj_5249, n135_adj_5250, 
        n138_adj_5251, n141_adj_5252, n144_adj_5253, n147_adj_5254, 
        n150_adj_5255, n153_adj_5256, n156_adj_5257, n159_adj_5258, 
        n162_adj_5259, n165_adj_5260, n168_adj_5261, n171_adj_5262, 
        n174_adj_5263, n177_adj_5264, n180_adj_5265, n183_adj_5266, 
        n78_adj_5267, n81_adj_5268, n84_adj_5269, n87_adj_5270, n90_adj_5271, 
        n93_adj_5272, n96_adj_5273, n99_adj_5274, n102_adj_5275, n105_adj_5276, 
        n108_adj_5277, n111_adj_5278, n114_adj_5279, n117_adj_5280, 
        n120_adj_5281, n123_adj_5282, n126_adj_5283, n129_adj_5284, 
        n132_adj_5285, n135_adj_5286, n138_adj_5287, n141_adj_5288, 
        n144_adj_5289, n147_adj_5290, n150_adj_5291, n153_adj_5292, 
        n156_adj_5293, n159_adj_5294, n162_adj_5295, n165_adj_5296, 
        n168_adj_5297, n171_adj_5298, n174_adj_5299, n177_adj_5300, 
        n180_adj_5301, n183_adj_5302, cout_adj_5303, n16598, n16640, 
        n16597, n16639, n16596, n16411, n51_adj_5304, n54_adj_5305, 
        n16638, n57_adj_5306, n16595, n60_adj_5307, n63_adj_5308, 
        n16557, n66_adj_5309, n16637, n69_adj_5310, n72_adj_5311, 
        n75_adj_5312, n78_adj_5313, n81_adj_5314, n16636, n84_adj_5315, 
        n87_adj_5316, n90_adj_5317, n16339, n16635, n16594, n16593, 
        n16634, n16592, n16633, n16591, n16632, n12136, n16420, 
        n16590, n16410, n16589, n16573, n16588, n16484, n16483, 
        n16482, n16481, n16480, n16479, n16409, n16408, n16478, 
        n16477, n16407, n16587, n78_adj_5318, n16572, n81_adj_5319, 
        n84_adj_5320, n87_adj_5321, n90_adj_5322, n16474, n93_adj_5323, 
        n96_adj_5324, n99_adj_5325, n102_adj_5326, n17310, n105_adj_5327, 
        n16406, n108_adj_5328, n111_adj_5329, n16473, n114_adj_5330, 
        n117_adj_5331, n16472, n120_adj_5332, n123_adj_5333, n16405, 
        n126_adj_5334, n129_adj_5335, n16471, n132_adj_5336, n135_adj_5337, 
        n16470, n138_adj_5338, n141_adj_5339, n16586, n144_adj_5340, 
        n16571, n147_adj_5341, n150_adj_5342, n153_adj_5343, n156_adj_5344, 
        n159_adj_5345, n162_adj_5346, n165_adj_5347, n168_adj_5348, 
        n16585, n171_adj_5349, n174_adj_5350, n12059, n177_adj_5351, 
        n12057, n180_adj_5352, n12055, n183_adj_5353, n12049, n12047, 
        n16337, n12043, n12037, n12035, n12033, n12031, n12029, 
        n12025, n12023, n12021, n12019, n12017, n12015, n12013, 
        n12011, n12009, n12007, n12003, n12001, n11999, n11995, 
        n11993, n11989, n11985, n18129, n11981, n12223, n11973, 
        n11971, n11969, clk_80mhz_enable_891, n11965, n11963, n16584, 
        n16583, n78_adj_5354, n81_adj_5355, n84_adj_5356, n87_adj_5357, 
        n90_adj_5358, n93_adj_5359, n96_adj_5360, n99_adj_5361, n102_adj_5362, 
        n105_adj_5363, n108_adj_5364, n111_adj_5365, n114_adj_5366, 
        n117_adj_5367, n120_adj_5368, n123_adj_5369, n126_adj_5370, 
        n129_adj_5371, n132_adj_5372, n135_adj_5373, n138_adj_5374, 
        n141_adj_5375, n144_adj_5376, n147_adj_5377, n150_adj_5378, 
        n153_adj_5379, n156_adj_5380, n159_adj_5381, n162_adj_5382, 
        n165_adj_5383, n168_adj_5384, n171_adj_5385, n174_adj_5386, 
        n177_adj_5387, n180_adj_5388, n183_adj_5389, n130_adj_5390, 
        n133_adj_5391, n136_adj_5392, n139_adj_5393, n142_adj_5394, 
        n145_adj_5395, n148_adj_5396, n151_adj_5397, n154_adj_5398, 
        n157_adj_5399, n160_adj_5400, n163_adj_5401, n166_adj_5402, 
        n169_adj_5403, n16469, n172_adj_5404, n16468, n175_adj_5405, 
        n16467, n178_adj_5406, n16466, n181_adj_5407, n16465, n184_adj_5408, 
        n16464, n187_adj_5409, n16463, n190_adj_5410, n16462, n193_adj_5411, 
        n16461, n196_adj_5412, n16460, n199_adj_5413, n16459, n202_adj_5414, 
        n16458, n205_adj_5415, n16457, n208_adj_5416, n211_adj_5417, 
        n16630, n214_adj_5418, n16629, n217_adj_5419, n220_adj_5420, 
        n223_adj_5421, n16369, n226_adj_5422, n229_adj_5423, n232_adj_5424, 
        n235_adj_5425, n238_adj_5426, n241_adj_5427, n244_adj_5428, 
        n247_adj_5429, n250_adj_5430, n253_adj_5431, n256_adj_5432, 
        n259_adj_5433, n16563, n262_adj_5434, n265_adj_5435, n16453, 
        n268_adj_5436, n271_adj_5437, n16628, n274_adj_5438, n16627, 
        n277_adj_5439, n280_adj_5440, n283_adj_5441, n16562, n286_adj_5442, 
        n289_adj_5443, n292_adj_5444, n16626, n295_adj_5445, n16625, 
        n298_adj_5446, n16889, n301_adj_5447, n16452, n304, n16561, 
        n307, n16888, n310, n16624, n313, n16623, n316, n16570, 
        n16887, n16622, n16582, n16886, n16885, n16621, n16404, 
        n16620, n16884, n11716, n16619, n16618, n16883, n16351, 
        n16617, n16569, n16403, n16882, n16616, n16615, n16451, 
        n16881, n16450, n15420, n16560, n16559, n16402, n16614, 
        n16613, n16612, n16611, n16558, n16875, n16216, n16215, 
        n16214, n16213, n16212, n16211, n16210, n16209, n16208, 
        n16207, n16206, n16205, n16204, n16203, n16202, n16201, 
        n78_adj_5448, n81_adj_5449, n84_adj_5450, n87_adj_5451, n90_adj_5452, 
        n93_adj_5453, n96_adj_5454, n99_adj_5455, n102_adj_5456, n105_adj_5457, 
        n108_adj_5458, n111_adj_5459, n114_adj_5460, n16874, n117_adj_5461, 
        n120_adj_5462, n16873, n123_adj_5463, n16610, n126_adj_5464, 
        n16449, n129_adj_5465, n16448, n132_adj_5466, n135_adj_5467, 
        n16872, n138_adj_5468, n141_adj_5469, n16401, n144_adj_5470, 
        n147_adj_5471, n16871, n150_adj_5472, n16870, n153_adj_5473, 
        n16609, n156_adj_5474, n16400, n159_adj_5475, n16608, n162_adj_5476, 
        n16869, n165_adj_5477, n16868, n168_adj_5478, n171_adj_5479, 
        n174_adj_5480, n177_adj_5481, n16867, n180_adj_5482, n183_adj_5483, 
        n16447, n16607, n16606, n16446, n16399, n16568, n16605, 
        n16604, n16373, n16445, n16603, clk_80mhz_enable_831, n16861, 
        n16398, n16382, n16444, n16443, n16442, n16441, n16440, 
        n16439, n16438, n16437, n16436, n16433, n16432, n16431, 
        n16430, n16860, n16859, n16429, n16602, n16601, n16397, 
        n16858, n16857, n16600, n16428, n16427, n16426, n16425, 
        n16424, n16423, n16422, n16421, n16390, n16396, n11_adj_5484, 
        n44, n13_adj_5485, n47, n50, n16567, n53, n16581, n56, 
        n59, n62, n16856, n65_adj_5486, n16855, n16854, n16853, 
        n16580, n16370, n16847, n16846, n16845, n16844, n16843, 
        n16842, n16841, n16395, n16840, n16566, n16579, n16578, 
        n16834, n16565, n16833, n16394, n11_adj_5487, n16832, n13_adj_5488, 
        n16831, n16577, n16830, n16393, n16829, n16828, n18145, 
        n16392, n16822, n16821, n16820, n16200, n16819, n16818, 
        n16817, n16816, n16199, n16815, n16198, n16813, n16812, 
        n16811, n16810, n16809, n16808, n16807, n12912, n16806, 
        n16805, n16799, n16576, n16798, n16797, n16796, n16575, 
        n16197, n16196, n16195, n16194, n16193, n16192, n16191, 
        n16190, n16189, n16188, n16187, n16186, n16185, n16184, 
        n16183, n16182, n16181, n16180, n16179, n16178, n16177, 
        n16176, n16175, n16174, n16173, n16172, n16171, n16170, 
        n16169, n16168, n16167, n16166, n16165, n16164, n16163, 
        n16162, n16161, n16160, n16159, n16158, n16157, n16156, 
        n16155, n16154, n16153, n16152, n16151, n16150, n16149, 
        n16148, n16147, n16146, n16145, n16144, n16143, n16142, 
        n16141, n16140, n16139, n16138, n16137, n16136, n16135, 
        n16134, n16133, n16132, n16131, n16130, n16129, n16128, 
        n16127, n16126, n16125, n16124, n16123, n16122, n16121, 
        n16120, n16119, n16118, n16117, n16116, n16115, n16114, 
        n16113, n16112, n16111, n16110, n16109, n16108, n16107, 
        n16106, n16105, n16104, n16103, n16102, n16101, n16100, 
        n16099, n16098, n16097, n16096, n16095, n16094, n16093, 
        n16092, n16091, n16090, n16089, n16088, n16087, n16086, 
        n16085, n16084, n16083, n16082, n16081, n16080, n16079, 
        n16078, n16077, n16076, n16075, n16074, n16073, n16072, 
        n16071, n16070, n16069, n16068, n16067, n16066, n16065, 
        n16064, n16063, n16062, n16061, n16060, n16059, n16058, 
        n16057, n16056, n16053, n16052, n16051, n16050, n16049, 
        n16048, n16047, n16046, n16045, n16044, n16043, n16042, 
        n16041, n16040, n16039, n16038, n16037, n16036, n16031, 
        n16030, n16029, n16028, n16027, n16026, n16025, n16024, 
        n16023, n16022, n16021, n16020, n16019, n16018, n16017, 
        n16016, n16015, n16014, n16010, n16009, n16008, n16007, 
        n16006, n16005, n16004, n16003, n16002, n16001, n16000, 
        n15999, n15998, n15997, n15996, n15995, n15994, n15993, 
        n15992, n15991, n15990, n15989, n15988, n15987, n15986, 
        n15985, n15984, n15983, n15982, n15981, n15980, n15979, 
        n15978, n15977, n15976, n15975, n15974, n15973, n15972, 
        n15971, n15970, n15969, n15968, n15967, n15966, n15965, 
        n15964, n15963, n15962, n15961, n15960, n15959, n15958, 
        n15957, cout_adj_5489, n15955, n15954, n15953, n15952, n15951, 
        n15950, n15949, n15948, n15947, n15946, n15945, n15944, 
        n15943, n15942, n15941, n15940, n15939, n15938, n15934, 
        n15933, n15932, n15931, n15930, n15929, n15928, n15927, 
        n15926, n15925, n15924, n15923, n15922, n15921, n15920, 
        n15919, n15918, n15917, n15916, n15915, n15914, n15913, 
        n15912, n15911, n15910, n15909, n15908, n15907, n15906, 
        n15905, n15904, n15903, n15902, n15901, n15900, n15899, 
        n15897, n15896, n15895, n15894, n15893, n15892, n15891, 
        n15890, n15889, n15888, n15887, n15886, n15885, n15884, 
        n15883, n15882, n15881, n15880, n15876, n15875, n15874, 
        n15873, n15872, n15871, n15870, n15869, n15868, n15867, 
        n15866, n15865, n15864, n15863, n15862, n15861, n15860, 
        n15859, n15857, n15856, n15855, n15854, n15853, n15852, 
        n15851, n15850, n15849, n15848, n15847, n15846, n15845, 
        n15844, n15843, cout_adj_5490, n15842, n15841, n15840, n15835, 
        n15834, n15833, n15832, n15831, n15830, n15829, n15828, 
        n15827, n15826, n15825, n15824, n15823, n15822, n15821, 
        n15820, n15819, n15818, n15814, n15813, n15812, n15811, 
        n15810, n15809, n15808, n15807, n15806, n15805, n15804, 
        n15803, n15802, n15801, n15800, n15799, n15798, n15797, 
        n15796, n15795, n52, n15794, n55, n15793, n58, n15792, 
        n61, n15791, n64_adj_5491, n15790, n67, n15789, n70, n15788, 
        n73, n15787, n76_adj_5492, n15786, n79_adj_5493, n15785, 
        n82_adj_5494, n15784, n85_adj_5495, n15783, n15782, n15781, 
        n15780, n15779, n15778, n15777, n15776, n15775, n15774, 
        n15773, n15772, n15771, n15770, n15769, n15768, n15767, 
        n15766, n15765, n15764, n15763, n15762, n15761, n15759, 
        n15758, n15757, n15756, n15755, n15754, n15753, n15752, 
        n15751, n15750, n15749, n15748, n15747, n15746, n15745, 
        n15744, n15743, n15742, n15738, n15737, n15736, n15735, 
        n15734, n15733, n15732, n15731, n15730, n15729, n15728, 
        n15727, n15726, n15725, n15724, n15723, n15722, n15721, 
        n15720, n15719, n15718, n15717, n15716, n15715, n15714, 
        n15713, n15712, n15711, n15710, n15709, n15708, n15707, 
        n15706, n15705, n15704, n15703, n15701, n15700, n15699, 
        n15698, n15697, n15696, n15695, n15694, n15693, n15692, 
        n15691, n15690, n15689, n15688, n15687, n15686, n15685, 
        cout_adj_5496, n15684, n15680, n15679, n15678, n15677, n15676, 
        n15675, n15674, n15673, n15672, n15671, n15670, n15669, 
        n15668, n15667, n15666, n15665, n15664, n15663, n15661, 
        n15660, n15659, n15658, n15657, n15656, n15655, n15654, 
        n15653, n15652, n15651, n15650, n15649, n15648, n15647, 
        n15646, n15645, n15644, n15642, n15641, n15640, n15639, 
        n15638, n15637, n15636, n15635, n15634, n15633, n45_adj_5497, 
        n15632, n48_adj_5498, n15631, n51_adj_5499, n15630, n54_adj_5500, 
        n15629, n57_adj_5501, n15628, n60_adj_5502, n15627, n63_adj_5503, 
        n15626, n66_adj_5504, n15625, n69_adj_5505, n15624, n72_adj_5506, 
        n15623, n75_adj_5507, n15622, n78_adj_5508, n15621, n81_adj_5509, 
        n15620, n84_adj_5510, n15619, n87_adj_5511, n15618, n90_adj_5512, 
        n15617, n15616, n15615, n15614, n15613, n15612, n15611, 
        n15610, n15609, n15608, n15607, n15606, n15605, n15604, 
        n15603, n15602, n15601, n15600, n15599, n15597, n15596, 
        n15595, n15594, n15593, n15592, n15591, n15590, n15589, 
        n15588, n15587, n15586, n15585, n15584, n15583, n15582, 
        n15581, n15580, n15579, n15578, n15577, n15576, n15575, 
        n45_adj_5513, n48_adj_5514, n15574, n51_adj_5515, n15573, 
        n54_adj_5516, n15572, n57_adj_5517, n15571, n60_adj_5518, 
        n15570, n63_adj_5519, n15569, n66_adj_5520, n15568, n69_adj_5521, 
        n15567, n72_adj_5522, n15566, n75_adj_5523, n15565, n78_adj_5524, 
        n15564, n81_adj_5525, n15563, n84_adj_5526, n15562, n87_adj_5527, 
        n15560, n90_adj_5528, n15559, n15558, n15557, n15556, n15555, 
        n15554, n15553, n15552, n15551, n15550, n15549, n15548, 
        n15547, n15546, n15545, n15544, n15543, n15541, n15540, 
        n15539, n15538, n15537, n15536, n15535, n15534, n15533, 
        n15532, n15531, n15530, n15529, n15528, n15527, n15526, 
        n15525, n15524, n45_adj_5529, n48_adj_5530, n15520, n51_adj_5531, 
        n15519, n54_adj_5532, n15518, n57_adj_5533, n15517, n60_adj_5534, 
        n15516, n63_adj_5535, n15515, n66_adj_5536, n15514, n69_adj_5537, 
        n15513, n72_adj_5538, n15512, n75_adj_5539, n15511, n78_adj_5540, 
        n15510, n81_adj_5541, n15509, n84_adj_5542, n15508, n87_adj_5543, 
        n15507, n90_adj_5544, n15506, n15505, n15504, n15503, n15501, 
        n15500, n15499, n15498, n15497, n15496, n15495, n15494, 
        n15493, n15492, n15491, n15490, n15489, n15488, n15487, 
        n15486, n15485, n15484, n15483, n15482, n15481, n15480, 
        n15479, n15478, n15477, n15476, n15475, n15474, n15473, 
        n15472, n15471, n15470, n15469, n15468, n15467, n15466, 
        n15465, n15464, n15463, n15462, n15461, n15460, n15459, 
        n15458, n15457, n15456, n15455, n15454, n15453, n15452, 
        n15451, n15450, n15449, n15448, n15447, n15446, n15445, 
        n15444, n15443, n15442, n15441, n15440, n15439, n15438, 
        n15437, n15436, n15435, n15434, n15433, n15432, n15431, 
        n15430, n15429, n15428, n15427, n15426, n15425, n15424, 
        n15423, n15422, n15421, n18087, n18086, n76_adj_5545, n79_adj_5546, 
        n82_adj_5547, n85_adj_5548, n88_adj_5549, n91_adj_5550, n94_adj_5551, 
        n97_adj_5552, n100_adj_5553, n103_adj_5554, n106_adj_5555, n109_adj_5556, 
        n112_adj_5557, n115_adj_5558, n118_adj_5559, n17536, n17595, 
        n17593, n45_adj_5560, n48_adj_5561, n51_adj_5562, n18075, 
        n54_adj_5563, n57_adj_5564, n60_adj_5565, n63_adj_5566, n66_adj_5567, 
        n69_adj_5568, n72_adj_5569, n75_adj_5570, n78_adj_5571, n81_adj_5572, 
        n84_adj_5573, n87_adj_5574, n90_adj_5575, n18074, n78_adj_5576, 
        n81_adj_5577, n84_adj_5578, n87_adj_5579, n90_adj_5580, n93_adj_5581, 
        n96_adj_5582, n99_adj_5583, n102_adj_5584, n105_adj_5585, n108_adj_5586, 
        n111_adj_5587, n114_adj_5588, n117_adj_5589, n120_adj_5590, 
        n123_adj_5591, n126_adj_5592, n129_adj_5593, n132_adj_5594, 
        n135_adj_5595, n138_adj_5596, n141_adj_5597, n144_adj_5598, 
        n147_adj_5599, n150_adj_5600, n153_adj_5601, n156_adj_5602, 
        n159_adj_5603, n162_adj_5604, n165_adj_5605, n168_adj_5606, 
        n171_adj_5607, n174_adj_5608, n177_adj_5609, n180_adj_5610, 
        n183_adj_5611, n15419, n15418, n15417, n18144, n18143, n15416, 
        n15415, n15414, n15413, n15412, n17805, n15409, n15408, 
        n15407, cout_adj_5612, n15406, n15405, n15404, n15403, n15402, 
        n15400, n15395, n48_adj_5613, n51_adj_5614, n54_adj_5615, 
        n57_adj_5616, n60_adj_5617, n63_adj_5618, n66_adj_5619, n69_adj_5620, 
        n72_adj_5621, n75_adj_5622, n15394, n15364, n15397, n78_adj_5623, 
        n81_adj_5624, n84_adj_5625, n87_adj_5626, n90_adj_5627, n93_adj_5628, 
        n96_adj_5629, n99_adj_5630, n102_adj_5631, n105_adj_5632, n108_adj_5633, 
        n111_adj_5634, n114_adj_5635, n117_adj_5636, n120_adj_5637, 
        n123_adj_5638, n126_adj_5639, n129_adj_5640, n132_adj_5641, 
        n135_adj_5642, n138_adj_5643, n141_adj_5644, n144_adj_5645, 
        n147_adj_5646, n150_adj_5647, n153_adj_5648, n156_adj_5649, 
        n159_adj_5650, n162_adj_5651, n165_adj_5652, n168_adj_5653, 
        n171_adj_5654, n174_adj_5655, n177_adj_5656, n180_adj_5657, 
        n183_adj_5658, n15398, n18131, n15393, n15392, n17784, clk_80mhz_enable_1471, 
        clk_80mhz_enable_881, n18127, n18142, n17496, n26_adj_5659, 
        n7_adj_5660, n15401, n8_adj_5661, n15399, n10_adj_5662, n15396, 
        n18301, n18141, clk_80mhz_enable_1470, n18268, n17298, n18139, 
        n18138, cout_adj_5663, n13099;
    
    VHI i2 (.Z(VCC_net));
    Mixer Mixer1 (.MixerOutSin({MixerOutSin}), .clk_80mhz(clk_80mhz), .DiffOut_c(DiffOut_c), 
          .MixerOutCos({MixerOutCos}), .RFIn_c(RFIn_c), .\LOSine[2] (LOSine[2]), 
          .MixerOutSin_11__N_236({MixerOutSin_11__N_236}), .\LOSine[3] (LOSine[3]), 
          .\LOSine[4] (LOSine[4]), .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), 
          .\LOSine[7] (LOSine[7]), .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), 
          .\LOSine[10] (LOSine[10]), .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), 
          .\LOCosine[2] (LOCosine[2]), .MixerOutCos_11__N_250({MixerOutCos_11__N_250}), 
          .\LOCosine[3] (LOCosine[3]), .\LOCosine[1] (LOCosine[1]), .\LOCosine[4] (LOCosine[4]), 
          .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
          .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
          .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
          .\LOSine[1] (LOSine[1])) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(170[7] 178[2])
    CCU2C _add_1_1439_add_4_4 (.A0(d4_adj_5676[2]), .B0(d3_adj_5675[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[3]), .B1(d3_adj_5675[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16477), .COUT(n16478), .S0(d4_71__N_634_adj_5692[2]), 
          .S1(d4_71__N_634_adj_5692[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_2 (.A0(d4_adj_5676[0]), .B0(d3_adj_5675[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[1]), .B1(d3_adj_5675[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16477), .S1(d4_71__N_634_adj_5692[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1439_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_21 (.A0(d7[54]), .B0(cout_adj_5050), .C0(n129_adj_4941), 
          .D0(n19_adj_4569), .A1(d7[55]), .B1(cout_adj_5050), .C1(n126_adj_4940), 
          .D1(n18_adj_4570), .CIN(n16425), .COUT(n16426), .S0(d8_71__N_1603[54]), 
          .S1(d8_71__N_1603[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_34 (.A0(d_d9_adj_5685[67]), .B0(d9_adj_5684[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[68]), .B1(d9_adj_5684[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16510), .COUT(n16511), .S0(n90_adj_4913), 
          .S1(n87_adj_4912));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_34.INJECT1_1 = "NO";
    CCU2C add_4107_5 (.A0(phase_inc_carrGen[2]), .B0(n13099), .C0(n2390), 
          .D0(n11716), .A1(phase_inc_carrGen[3]), .B1(n13099), .C1(n2389), 
          .D1(n11716), .CIN(n16720), .COUT(n16721), .S0(n317), .S1(n314));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_5.INIT0 = 16'h74b8;
    defparam add_4107_5.INIT1 = 16'h74b8;
    defparam add_4107_5.INJECT1_0 = "NO";
    defparam add_4107_5.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_10 (.A0(d4_adj_5676[43]), .B0(d3_adj_5675[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[44]), .B1(d3_adj_5675[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16271), .COUT(n16272), .S0(n162_adj_4558), 
          .S1(n159_adj_4559));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_7 (.A0(d_tmp_adj_5671[40]), .B0(cout_adj_5489), 
          .C0(n171_adj_5349), .D0(n33), .A1(d_tmp_adj_5671[41]), .B1(cout_adj_5489), 
          .C1(n168_adj_5348), .D1(n32), .CIN(n16459), .COUT(n16460), 
          .S0(d6_71__N_1459_adj_5705[40]), .S1(d6_71__N_1459_adj_5705[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_23 (.A0(d_tmp[56]), .B0(cout_adj_5496), .C0(n123_adj_5066), 
          .D0(n17_adj_4732), .A1(d_tmp[57]), .B1(cout_adj_5496), .C1(n120_adj_5065), 
          .D1(n16_adj_4731), .CIN(n16334), .COUT(n16335), .S0(d6_71__N_1459[56]), 
          .S1(d6_71__N_1459[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_5 (.A0(d_tmp_adj_5671[38]), .B0(cout_adj_5489), 
          .C0(n177_adj_5351), .D0(n35), .A1(d_tmp_adj_5671[39]), .B1(cout_adj_5489), 
          .C1(n174_adj_5350), .D1(n34), .CIN(n16458), .COUT(n16459), 
          .S0(d6_71__N_1459_adj_5705[38]), .S1(d6_71__N_1459_adj_5705[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_5.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    CCU2C _add_1_1448_add_4_21 (.A0(d_tmp[54]), .B0(cout_adj_5496), .C0(n129_adj_5068), 
          .D0(n19_adj_4808), .A1(d_tmp[55]), .B1(cout_adj_5496), .C1(n126_adj_5067), 
          .D1(n18_adj_4809), .CIN(n16333), .COUT(n16334), .S0(d6_71__N_1459[54]), 
          .S1(d6_71__N_1459[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_21.INJECT1_1 = "NO";
    FD1S3AX o_Rx_DV_40 (.D(o_Rx_DV1), .CK(clk_80mhz), .Q(o_Rx_DV));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_DV_40.GSR = "ENABLED";
    CCU2C add_4107_3 (.A0(phase_inc_carrGen[0]), .B0(n13099), .C0(n17496), 
          .D0(n18131), .A1(phase_inc_carrGen[1]), .B1(n13099), .C1(n2391), 
          .D1(n3716), .CIN(n16719), .COUT(n16720), .S0(n323), .S1(n320));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_3.INIT0 = 16'h74b8;
    defparam add_4107_3.INIT1 = 16'h74b8;
    defparam add_4107_3.INJECT1_0 = "NO";
    defparam add_4107_3.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16494), .S0(cout_adj_5149));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1439_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1439_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_19 (.A0(d7[52]), .B0(cout_adj_5050), .C0(n135_adj_4943), 
          .D0(n21_adj_4567), .A1(d7[53]), .B1(cout_adj_5050), .C1(n132_adj_4942), 
          .D1(n20_adj_4568), .CIN(n16424), .COUT(n16425), .S0(d8_71__N_1603[52]), 
          .S1(d8_71__N_1603[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_36 (.A0(d4_adj_5676[34]), .B0(d3_adj_5675[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[35]), .B1(d3_adj_5675[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16493), .COUT(n16494), .S0(d4_71__N_634_adj_5692[34]), 
          .S1(d4_71__N_634_adj_5692[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_34 (.A0(d4_adj_5676[32]), .B0(d3_adj_5675[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[33]), .B1(d3_adj_5675[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16492), .COUT(n16493), .S0(d4_71__N_634_adj_5692[32]), 
          .S1(d4_71__N_634_adj_5692[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_34.INJECT1_1 = "NO";
    LUT4 mux_326_i29_4_lut (.A(n12003), .B(n235_adj_5425), .C(n18135), 
         .D(n2593), .Z(n2364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i29_4_lut.init = 16'hcfca;
    CCU2C _add_1_1439_add_4_30 (.A0(d4_adj_5676[28]), .B0(d3_adj_5675[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[29]), .B1(d3_adj_5675[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16490), .COUT(n16491), .S0(d4_71__N_634_adj_5692[28]), 
          .S1(d4_71__N_634_adj_5692[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5489), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16457));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1481_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1481_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_1.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[54]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    CCU2C _add_1_1442_add_4_32 (.A0(d5_adj_5677[30]), .B0(d4_adj_5676[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[31]), .B1(d4_adj_5676[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16450), .COUT(n16451), .S0(d5_71__N_706_adj_5693[30]), 
          .S1(d5_71__N_706_adj_5693[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_32.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[52]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    CCU2C _add_1_1442_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16453), .S0(cout_adj_5150));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1442_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1442_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_cout.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    CCU2C _add_1_1442_add_4_26 (.A0(d5_adj_5677[24]), .B0(d4_adj_5676[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[25]), .B1(d4_adj_5676[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16447), .COUT(n16448), .S0(d5_71__N_706_adj_5693[24]), 
          .S1(d5_71__N_706_adj_5693[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_17 (.A0(d7[50]), .B0(cout_adj_5050), .C0(n141_adj_4945), 
          .D0(n23), .A1(d7[51]), .B1(cout_adj_5050), .C1(n138_adj_4944), 
          .D1(n22_adj_4836), .CIN(n16423), .COUT(n16424), .S0(d8_71__N_1603[50]), 
          .S1(d8_71__N_1603[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_17.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[50]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    PWM PWM1 (.\DemodOut[9] (DemodOut[9]), .\DataInReg[0] (DataInReg[0]), 
        .clk_80mhz(clk_80mhz), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
        .counter({counter}), .GND_net(GND_net), .VCC_net(VCC_net), .\DataInReg[1] (DataInReg[1]), 
        .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg[2] (DataInReg[2]), 
        .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg[3] (DataInReg[3]), 
        .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg[4] (DataInReg[4]), 
        .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg[5] (DataInReg[5]), 
        .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg[6] (DataInReg[6]), 
        .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg[7] (DataInReg[7]), 
        .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg[8] (DataInReg[8]), 
        .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DataInReg[9] (DataInReg[9])) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(199[5] 205[2])
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    CCU2C _add_1_1481_add_4_3 (.A0(d_tmp_adj_5671[36]), .B0(cout_adj_5489), 
          .C0(n183_adj_5353), .D0(n37), .A1(d_tmp_adj_5671[37]), .B1(cout_adj_5489), 
          .C1(n180_adj_5352), .D1(n36), .CIN(n16457), .COUT(n16458), 
          .S0(d6_71__N_1459_adj_5705[36]), .S1(d6_71__N_1459_adj_5705[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_3.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[48]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    CCU2C _add_1_1448_add_4_19 (.A0(d_tmp[52]), .B0(cout_adj_5496), .C0(n135_adj_5070), 
          .D0(n21_adj_4806), .A1(d_tmp[53]), .B1(cout_adj_5496), .C1(n132_adj_5069), 
          .D1(n20_adj_4807), .CIN(n16332), .COUT(n16333), .S0(d6_71__N_1459[52]), 
          .S1(d6_71__N_1459[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_34 (.A0(d5_adj_5677[32]), .B0(d4_adj_5676[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[33]), .B1(d4_adj_5676[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16451), .COUT(n16452), .S0(d5_71__N_706_adj_5693[32]), 
          .S1(d5_71__N_706_adj_5693[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_22 (.A0(d5_adj_5677[20]), .B0(d4_adj_5676[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[21]), .B1(d4_adj_5676[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16445), .COUT(n16446), .S0(d5_71__N_706_adj_5693[20]), 
          .S1(d5_71__N_706_adj_5693[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_36 (.A0(d5_adj_5677[34]), .B0(d4_adj_5676[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[35]), .B1(d4_adj_5676[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16452), .COUT(n16453), .S0(d5_71__N_706_adj_5693[34]), 
          .S1(d5_71__N_706_adj_5693[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_17 (.A0(d_tmp[50]), .B0(cout_adj_5496), .C0(n141_adj_5072), 
          .D0(n23_adj_4804), .A1(d_tmp[51]), .B1(cout_adj_5496), .C1(n138_adj_5071), 
          .D1(n22_adj_4805), .CIN(n16331), .COUT(n16332), .S0(d6_71__N_1459[50]), 
          .S1(d6_71__N_1459[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_28 (.A0(d4_adj_5676[61]), .B0(d3_adj_5675[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[62]), .B1(d3_adj_5675[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16280), .COUT(n16281), .S0(n108_adj_4591), 
          .S1(n105_adj_4590));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_8 (.A0(d4_adj_5676[41]), .B0(d3_adj_5675[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[42]), .B1(d3_adj_5675[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16270), .COUT(n16271), .S0(n168_adj_4556), 
          .S1(n165_adj_4557));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_8.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[46]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[44]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    CCU2C _add_1_1442_add_4_20 (.A0(d5_adj_5677[18]), .B0(d4_adj_5676[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[19]), .B1(d4_adj_5676[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16444), .COUT(n16445), .S0(d5_71__N_706_adj_5693[18]), 
          .S1(d5_71__N_706_adj_5693[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_30 (.A0(d5_adj_5677[28]), .B0(d4_adj_5676[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[29]), .B1(d4_adj_5676[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16449), .COUT(n16450), .S0(d5_71__N_706_adj_5693[28]), 
          .S1(d5_71__N_706_adj_5693[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_18 (.A0(d1_adj_5673[51]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[52]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16081), .COUT(n16082), .S0(n138_adj_5596), 
          .S1(n135_adj_5595));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_18.INJECT1_1 = "NO";
    LUT4 i2248_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(n18268), .D(n301), 
         .Z(n11963)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2248_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1442_add_4_28 (.A0(d5_adj_5677[26]), .B0(d4_adj_5676[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[27]), .B1(d4_adj_5676[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16448), .COUT(n16449), .S0(d5_71__N_706_adj_5693[26]), 
          .S1(d5_71__N_706_adj_5693[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_15 (.A0(d_tmp[48]), .B0(cout_adj_5496), .C0(n147_adj_5074), 
          .D0(n25_adj_4802), .A1(d_tmp[49]), .B1(cout_adj_5496), .C1(n144_adj_5073), 
          .D1(n24_adj_4803), .CIN(n16330), .COUT(n16331), .S0(d6_71__N_1459[48]), 
          .S1(d6_71__N_1459[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_16 (.A0(d1_adj_5673[49]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[50]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16080), .COUT(n16081), .S0(n144_adj_5598), 
          .S1(n141_adj_5597));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_16.INJECT1_1 = "NO";
    FD1P3AX CICGain__i1 (.D(led_c_0), .SP(clk_80mhz_enable_1470), .CK(clk_80mhz), 
            .Q(CICGain[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam CICGain__i1.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[42]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    CCU2C _add_1_1490_add_4_33 (.A0(d4_adj_5676[66]), .B0(cout_adj_5150), 
          .C0(n93_adj_4842), .D0(d5_adj_5677[66]), .A1(d4_adj_5676[67]), 
          .B1(cout_adj_5150), .C1(n90_adj_4841), .D1(d5_adj_5677[67]), 
          .CIN(n16361), .COUT(n16362), .S0(d5_71__N_706_adj_5693[66]), 
          .S1(d5_71__N_706_adj_5693[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_33.INJECT1_1 = "NO";
    LUT4 mux_326_i30_4_lut (.A(n2563), .B(n232_adj_5424), .C(n18135), 
         .D(n2593), .Z(n2363)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i30_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1568_add_4_14 (.A0(d1_adj_5673[47]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[48]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16079), .COUT(n16080), .S0(n150_adj_5600), 
          .S1(n147_adj_5599));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_32 (.A0(d4_adj_5676[30]), .B0(d3_adj_5675[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[31]), .B1(d3_adj_5675[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16491), .COUT(n16492), .S0(d4_71__N_634_adj_5692[30]), 
          .S1(d4_71__N_634_adj_5692[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_12 (.A0(d1_adj_5673[45]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[46]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16078), .COUT(n16079), .S0(n156_adj_5602), 
          .S1(n153_adj_5601));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_18 (.A0(d4_adj_5676[16]), .B0(d3_adj_5675[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[17]), .B1(d3_adj_5675[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16484), .COUT(n16485), .S0(d4_71__N_634_adj_5692[16]), 
          .S1(d4_71__N_634_adj_5692[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5150), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16346));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1490_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1490_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_16 (.A0(d4_adj_5676[14]), .B0(d3_adj_5675[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[15]), .B1(d3_adj_5675[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16483), .COUT(n16484), .S0(d4_71__N_634_adj_5692[14]), 
          .S1(d4_71__N_634_adj_5692[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_14 (.A0(d4_adj_5676[12]), .B0(d3_adj_5675[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[13]), .B1(d3_adj_5675[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16482), .COUT(n16483), .S0(d4_71__N_634_adj_5692[12]), 
          .S1(d4_71__N_634_adj_5692[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_12 (.A0(d4_adj_5676[10]), .B0(d3_adj_5675[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[11]), .B1(d3_adj_5675[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16481), .COUT(n16482), .S0(d4_71__N_634_adj_5692[10]), 
          .S1(d4_71__N_634_adj_5692[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_10 (.A0(d4_adj_5676[8]), .B0(d3_adj_5675[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[9]), .B1(d3_adj_5675[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16480), .COUT(n16481), .S0(d4_71__N_634_adj_5692[8]), 
          .S1(d4_71__N_634_adj_5692[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_24 (.A0(d5_adj_5677[22]), .B0(d4_adj_5676[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[23]), .B1(d4_adj_5676[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16446), .COUT(n16447), .S0(d5_71__N_706_adj_5693[22]), 
          .S1(d5_71__N_706_adj_5693[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_15 (.A0(d7[48]), .B0(cout_adj_5050), .C0(n147_adj_4947), 
          .D0(n25), .A1(d7[49]), .B1(cout_adj_5050), .C1(n144_adj_4946), 
          .D1(n24), .CIN(n16422), .COUT(n16423), .S0(d8_71__N_1603[48]), 
          .S1(d8_71__N_1603[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_31 (.A0(d4_adj_5676[64]), .B0(cout_adj_5150), 
          .C0(n99_adj_4844), .D0(d5_adj_5677[64]), .A1(d4_adj_5676[65]), 
          .B1(cout_adj_5150), .C1(n96_adj_4843), .D1(d5_adj_5677[65]), 
          .CIN(n16360), .COUT(n16361), .S0(d5_71__N_706_adj_5693[64]), 
          .S1(d5_71__N_706_adj_5693[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_13 (.A0(d_tmp[46]), .B0(cout_adj_5496), .C0(n153_adj_5076), 
          .D0(n27_adj_4800), .A1(d_tmp[47]), .B1(cout_adj_5496), .C1(n150_adj_5075), 
          .D1(n26_adj_4801), .CIN(n16329), .COUT(n16330), .S0(d6_71__N_1459[46]), 
          .S1(d6_71__N_1459[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_11 (.A0(d_tmp[44]), .B0(cout_adj_5496), .C0(n159_adj_5078), 
          .D0(n29_adj_4798), .A1(d_tmp[45]), .B1(cout_adj_5496), .C1(n156_adj_5077), 
          .D1(n28_adj_4799), .CIN(n16328), .COUT(n16329), .S0(d6_71__N_1459[44]), 
          .S1(d6_71__N_1459[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_11.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    CCU2C _add_1_1439_add_4_8 (.A0(d4_adj_5676[6]), .B0(d3_adj_5675[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[7]), .B1(d3_adj_5675[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16479), .COUT(n16480), .S0(d4_71__N_634_adj_5692[6]), 
          .S1(d4_71__N_634_adj_5692[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_6 (.A0(d4_adj_5676[4]), .B0(d3_adj_5675[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[5]), .B1(d3_adj_5675[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16478), .COUT(n16479), .S0(d4_71__N_634_adj_5692[4]), 
          .S1(d4_71__N_634_adj_5692[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_9 (.A0(d_tmp[42]), .B0(cout_adj_5496), .C0(n165_adj_5080), 
          .D0(n31_adj_4796), .A1(d_tmp[43]), .B1(cout_adj_5496), .C1(n162_adj_5079), 
          .D1(n30_adj_4797), .CIN(n16327), .COUT(n16328), .S0(d6_71__N_1459[42]), 
          .S1(d6_71__N_1459[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_9.INJECT1_1 = "NO";
    CCU2C add_4107_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n18127), .B1(n12912), .C1(led_c_4), .D1(n2845), .COUT(n16719));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_1.INIT0 = 16'h0000;
    defparam add_4107_1.INIT1 = 16'hf7ff;
    defparam add_4107_1.INJECT1_0 = "NO";
    defparam add_4107_1.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_7 (.A0(d_tmp[40]), .B0(cout_adj_5496), .C0(n171_adj_5082), 
          .D0(n33_adj_4794), .A1(d_tmp[41]), .B1(cout_adj_5496), .C1(n168_adj_5081), 
          .D1(n32_adj_4795), .CIN(n16326), .COUT(n16327), .S0(d6_71__N_1459[40]), 
          .S1(d6_71__N_1459[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_11 (.A0(d_tmp_adj_5671[44]), .B0(cout_adj_5489), 
          .C0(n159_adj_5345), .D0(n29_adj_2749), .A1(d_tmp_adj_5671[45]), 
          .B1(cout_adj_5489), .C1(n156_adj_5344), .D1(n28_adj_2750), .CIN(n16461), 
          .COUT(n16462), .S0(d6_71__N_1459_adj_5705[44]), .S1(d6_71__N_1459_adj_5705[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_31 (.A0(d_tmp_adj_5671[64]), .B0(cout_adj_5489), 
          .C0(n99_adj_5325), .D0(n9), .A1(d_tmp_adj_5671[65]), .B1(cout_adj_5489), 
          .C1(n96_adj_5324), .D1(n8), .CIN(n16471), .COUT(n16472), .S0(d6_71__N_1459_adj_5705[64]), 
          .S1(d6_71__N_1459_adj_5705[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_5 (.A0(d_tmp[38]), .B0(cout_adj_5496), .C0(n177_adj_5084), 
          .D0(n35_adj_4810), .A1(d_tmp[39]), .B1(cout_adj_5496), .C1(n174_adj_5083), 
          .D1(n34_adj_4793), .CIN(n16325), .COUT(n16326), .S0(d6_71__N_1459[38]), 
          .S1(d6_71__N_1459[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_3 (.A0(d_tmp[36]), .B0(cout_adj_5496), .C0(n183_adj_5086), 
          .D0(n37_adj_4812), .A1(d_tmp[37]), .B1(cout_adj_5496), .C1(n180_adj_5085), 
          .D1(n36_adj_4811), .CIN(n16324), .COUT(n16325), .S0(d6_71__N_1459[36]), 
          .S1(d6_71__N_1459[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_3.INJECT1_1 = "NO";
    LUT4 i2344_3_lut_4_lut (.A(n18267), .B(n18138), .C(n18268), .D(n133), 
         .Z(n12059)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2344_3_lut_4_lut.init = 16'hfb0b;
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[40]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    CCU2C _add_1_1568_add_4_10 (.A0(d1_adj_5673[43]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[44]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16077), .COUT(n16078), .S0(n162_adj_5604), 
          .S1(n159_adj_5603));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_13 (.A0(d7[46]), .B0(cout_adj_5050), .C0(n153_adj_4949), 
          .D0(n27), .A1(d7[47]), .B1(cout_adj_5050), .C1(n150_adj_4948), 
          .D1(n26), .CIN(n16421), .COUT(n16422), .S0(d8_71__N_1603[46]), 
          .S1(d8_71__N_1603[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_18 (.A0(d5_adj_5677[16]), .B0(d4_adj_5676[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[17]), .B1(d4_adj_5676[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16443), .COUT(n16444), .S0(d5_71__N_706_adj_5693[16]), 
          .S1(d5_71__N_706_adj_5693[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5496), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16324));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1448_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1448_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_16 (.A0(d5_adj_5677[14]), .B0(d4_adj_5676[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[15]), .B1(d4_adj_5676[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16442), .COUT(n16443), .S0(d5_71__N_706_adj_5693[14]), 
          .S1(d5_71__N_706_adj_5693[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_10 (.A0(d5_adj_5677[8]), .B0(d4_adj_5676[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[9]), .B1(d4_adj_5676[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16439), .COUT(n16440), .S0(d5_71__N_706_adj_5693[8]), 
          .S1(d5_71__N_706_adj_5693[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_4 (.A0(d5_adj_5677[2]), .B0(d4_adj_5676[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[3]), .B1(d4_adj_5676[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16436), .COUT(n16437), .S0(d5_71__N_706_adj_5693[2]), 
          .S1(d5_71__N_706_adj_5693[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_11 (.A0(d7[44]), .B0(cout_adj_5050), .C0(n159_adj_4951), 
          .D0(n29), .A1(d7[45]), .B1(cout_adj_5050), .C1(n156_adj_4950), 
          .D1(n28), .CIN(n16420), .COUT(n16421), .S0(d8_71__N_1603[44]), 
          .S1(d8_71__N_1603[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_8 (.A0(d5_adj_5677[6]), .B0(d4_adj_5676[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[7]), .B1(d4_adj_5676[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16438), .COUT(n16439), .S0(d5_71__N_706_adj_5693[6]), 
          .S1(d5_71__N_706_adj_5693[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_14 (.A0(d5_adj_5677[12]), .B0(d4_adj_5676[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[13]), .B1(d4_adj_5676[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16441), .COUT(n16442), .S0(d5_71__N_706_adj_5693[12]), 
          .S1(d5_71__N_706_adj_5693[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_6 (.A0(d5_adj_5677[4]), .B0(d4_adj_5676[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[5]), .B1(d4_adj_5676[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16437), .COUT(n16438), .S0(d5_71__N_706_adj_5693[4]), 
          .S1(d5_71__N_706_adj_5693[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_2 (.A0(d5_adj_5677[0]), .B0(d4_adj_5676[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[1]), .B1(d4_adj_5676[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16436), .S1(d5_71__N_706_adj_5693[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1442_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_12 (.A0(d5_adj_5677[10]), .B0(d4_adj_5676[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[11]), .B1(d4_adj_5676[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16440), .COUT(n16441), .S0(d5_71__N_706_adj_5693[10]), 
          .S1(d5_71__N_706_adj_5693[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_8 (.A0(d1_adj_5673[41]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[42]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16076), .COUT(n16077), .S0(n168_adj_5606), 
          .S1(n165_adj_5605));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_9 (.A0(d7[42]), .B0(cout_adj_5050), .C0(n165_adj_4953), 
          .D0(n31_adj_4813), .A1(d7[43]), .B1(cout_adj_5050), .C1(n162_adj_4952), 
          .D1(n30), .CIN(n16419), .COUT(n16420), .S0(d8_71__N_1603[42]), 
          .S1(d8_71__N_1603[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_6 (.A0(d1_adj_5673[39]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[40]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16075), .COUT(n16076), .S0(n174_adj_5608), 
          .S1(n171_adj_5607));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_4 (.A0(d1_adj_5673[37]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[38]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16074), .COUT(n16075), .S0(n180_adj_5610), 
          .S1(n177_adj_5609));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_4.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(led_c_1), .B(led_c_4), .C(led_c_0), 
         .D(led_c_3), .Z(n17298)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2000;
    CCU2C _add_1_1568_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1_adj_5673[36]), .B1(MixerOutCos[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16074), .S1(n183_adj_5611));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1568_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16073), .S0(cout_adj_5087));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1421_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1421_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_cout.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    LUT4 mux_326_i27_4_lut (.A(n11999), .B(n241_adj_5427), .C(n18135), 
         .D(n2593), .Z(n2366)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i27_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1466_add_4_7 (.A0(d7[40]), .B0(cout_adj_5050), .C0(n171_adj_4955), 
          .D0(n33_adj_4696), .A1(d7[41]), .B1(cout_adj_5050), .C1(n168_adj_4954), 
          .D1(n32_adj_4792), .CIN(n16418), .COUT(n16419), .S0(d8_71__N_1603[40]), 
          .S1(d8_71__N_1603[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_29 (.A0(d4_adj_5676[62]), .B0(cout_adj_5150), 
          .C0(n105_adj_4846), .D0(d5_adj_5677[62]), .A1(d4_adj_5676[63]), 
          .B1(cout_adj_5150), .C1(n102_adj_4845), .D1(d5_adj_5677[63]), 
          .CIN(n16359), .COUT(n16360), .S0(d5_71__N_706_adj_5693[62]), 
          .S1(d5_71__N_706_adj_5693[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_5 (.A0(d7[38]), .B0(cout_adj_5050), .C0(n177_adj_4957), 
          .D0(n35_adj_4694), .A1(d7[39]), .B1(cout_adj_5050), .C1(n174_adj_4956), 
          .D1(n34_adj_4695), .CIN(n16417), .COUT(n16418), .S0(d8_71__N_1603[38]), 
          .S1(d8_71__N_1603[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_27 (.A0(d4_adj_5676[60]), .B0(cout_adj_5150), 
          .C0(n111_adj_4848), .D0(d5_adj_5677[60]), .A1(d4_adj_5676[61]), 
          .B1(cout_adj_5150), .C1(n108_adj_4847), .D1(d5_adj_5677[61]), 
          .CIN(n16358), .COUT(n16359), .S0(d5_71__N_706_adj_5693[60]), 
          .S1(d5_71__N_706_adj_5693[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_5 (.A0(d4_adj_5676[38]), .B0(cout_adj_5150), 
          .C0(n177_adj_4870), .D0(d5_adj_5677[38]), .A1(d4_adj_5676[39]), 
          .B1(cout_adj_5150), .C1(n174_adj_4869), .D1(d5_adj_5677[39]), 
          .CIN(n16347), .COUT(n16348), .S0(d5_71__N_706_adj_5693[38]), 
          .S1(d5_71__N_706_adj_5693[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_25 (.A0(d4_adj_5676[58]), .B0(cout_adj_5150), 
          .C0(n117_adj_4850), .D0(d5_adj_5677[58]), .A1(d4_adj_5676[59]), 
          .B1(cout_adj_5150), .C1(n114_adj_4849), .D1(d5_adj_5677[59]), 
          .CIN(n16357), .COUT(n16358), .S0(d5_71__N_706_adj_5693[58]), 
          .S1(d5_71__N_706_adj_5693[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_9 (.A0(d4_adj_5676[42]), .B0(cout_adj_5150), 
          .C0(n165_adj_4866), .D0(d5_adj_5677[42]), .A1(d4_adj_5676[43]), 
          .B1(cout_adj_5150), .C1(n162_adj_4865), .D1(d5_adj_5677[43]), 
          .CIN(n16349), .COUT(n16350), .S0(d5_71__N_706_adj_5693[42]), 
          .S1(d5_71__N_706_adj_5693[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_9.INJECT1_1 = "NO";
    LUT4 i2340_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(led_c_3), .D(n139), 
         .Z(n12055)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2340_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1466_add_4_37 (.A0(d7[70]), .B0(cout_adj_5050), .C0(n81_adj_4925), 
          .D0(n3_adj_4691), .A1(d7[71]), .B1(cout_adj_5050), .C1(n78_adj_4924), 
          .D1(n2_adj_4692), .CIN(n16433), .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_33 (.A0(d7[66]), .B0(cout_adj_5050), .C0(n93_adj_4929), 
          .D0(n7_adj_4658), .A1(d7[67]), .B1(cout_adj_5050), .C1(n90_adj_4928), 
          .D1(n6_adj_4687), .CIN(n16431), .COUT(n16432), .S0(d8_71__N_1603[66]), 
          .S1(d8_71__N_1603[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_31 (.A0(d7[64]), .B0(cout_adj_5050), .C0(n99_adj_4931), 
          .D0(n9_adj_4625), .A1(d7[65]), .B1(cout_adj_5050), .C1(n96_adj_4930), 
          .D1(n8_adj_4655), .CIN(n16430), .COUT(n16431), .S0(d8_71__N_1603[64]), 
          .S1(d8_71__N_1603[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_31.INJECT1_1 = "NO";
    LUT4 mux_326_i28_4_lut (.A(n12001), .B(n238_adj_5426), .C(n18135), 
         .D(n2593), .Z(n2365)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i28_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1421_add_4_36 (.A0(d4[34]), .B0(d3[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[35]), .B1(d3[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16072), .COUT(n16073), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_15 (.A0(d_tmp_adj_5671[48]), .B0(cout_adj_5489), 
          .C0(n147_adj_5341), .D0(n25_adj_2753), .A1(d_tmp_adj_5671[49]), 
          .B1(cout_adj_5489), .C1(n144_adj_5340), .D1(n24_adj_2754), .CIN(n16463), 
          .COUT(n16464), .S0(d6_71__N_1459_adj_5705[48]), .S1(d6_71__N_1459_adj_5705[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_37 (.A0(d3_adj_5675[70]), .B0(cout_adj_5149), 
          .C0(n81), .D0(d4_adj_5676[70]), .A1(d3_adj_5675[71]), .B1(cout_adj_5149), 
          .C1(n78), .D1(d4_adj_5676[71]), .CIN(n16319), .S0(d4_71__N_634_adj_5692[70]), 
          .S1(d4_71__N_634_adj_5692[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_35 (.A0(d3_adj_5675[68]), .B0(cout_adj_5149), 
          .C0(n87), .D0(d4_adj_5676[68]), .A1(d3_adj_5675[69]), .B1(cout_adj_5149), 
          .C1(n84), .D1(d4_adj_5676[69]), .CIN(n16318), .COUT(n16319), 
          .S0(d4_71__N_634_adj_5692[68]), .S1(d4_71__N_634_adj_5692[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_33 (.A0(d3_adj_5675[66]), .B0(cout_adj_5149), 
          .C0(n93), .D0(d4_adj_5676[66]), .A1(d3_adj_5675[67]), .B1(cout_adj_5149), 
          .C1(n90), .D1(d4_adj_5676[67]), .CIN(n16317), .COUT(n16318), 
          .S0(d4_71__N_634_adj_5692[66]), .S1(d4_71__N_634_adj_5692[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_31 (.A0(d3_adj_5675[64]), .B0(cout_adj_5149), 
          .C0(n99), .D0(d4_adj_5676[64]), .A1(d3_adj_5675[65]), .B1(cout_adj_5149), 
          .C1(n96), .D1(d4_adj_5676[65]), .CIN(n16316), .COUT(n16317), 
          .S0(d4_71__N_634_adj_5692[64]), .S1(d4_71__N_634_adj_5692[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_29 (.A0(d3_adj_5675[62]), .B0(cout_adj_5149), 
          .C0(n105_adj_4590), .D0(d4_adj_5676[62]), .A1(d3_adj_5675[63]), 
          .B1(cout_adj_5149), .C1(n102), .D1(d4_adj_5676[63]), .CIN(n16315), 
          .COUT(n16316), .S0(d4_71__N_634_adj_5692[62]), .S1(d4_71__N_634_adj_5692[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_37 (.A0(d_tmp_adj_5671[70]), .B0(cout_adj_5489), 
          .C0(n81_adj_5319), .D0(n3_adj_2760), .A1(d_tmp_adj_5671[71]), 
          .B1(cout_adj_5489), .C1(n78_adj_5318), .D1(n2_adj_2761), .CIN(n16474), 
          .S0(d6_71__N_1459_adj_5705[70]), .S1(d6_71__N_1459_adj_5705[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_34 (.A0(d4[32]), .B0(d3[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[33]), .B1(d3[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16071), .COUT(n16072), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_27 (.A0(d3_adj_5675[60]), .B0(cout_adj_5149), 
          .C0(n111_adj_4742), .D0(d4_adj_5676[60]), .A1(d3_adj_5675[61]), 
          .B1(cout_adj_5149), .C1(n108_adj_4591), .D1(d4_adj_5676[61]), 
          .CIN(n16314), .COUT(n16315), .S0(d4_71__N_634_adj_5692[60]), 
          .S1(d4_71__N_634_adj_5692[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_25 (.A0(d3_adj_5675[58]), .B0(cout_adj_5149), 
          .C0(n117_adj_4745), .D0(d4_adj_5676[58]), .A1(d3_adj_5675[59]), 
          .B1(cout_adj_5149), .C1(n114_adj_4744), .D1(d4_adj_5676[59]), 
          .CIN(n16313), .COUT(n16314), .S0(d4_71__N_634_adj_5692[58]), 
          .S1(d4_71__N_634_adj_5692[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_23 (.A0(d3_adj_5675[56]), .B0(cout_adj_5149), 
          .C0(n123_adj_4747), .D0(d4_adj_5676[56]), .A1(d3_adj_5675[57]), 
          .B1(cout_adj_5149), .C1(n120_adj_4746), .D1(d4_adj_5676[57]), 
          .CIN(n16312), .COUT(n16313), .S0(d4_71__N_634_adj_5692[56]), 
          .S1(d4_71__N_634_adj_5692[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_21 (.A0(d3_adj_5675[54]), .B0(cout_adj_5149), 
          .C0(n129_adj_4789), .D0(d4_adj_5676[54]), .A1(d3_adj_5675[55]), 
          .B1(cout_adj_5149), .C1(n126_adj_4788), .D1(d4_adj_5676[55]), 
          .CIN(n16311), .COUT(n16312), .S0(d4_71__N_634_adj_5692[54]), 
          .S1(d4_71__N_634_adj_5692[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_19 (.A0(d3_adj_5675[52]), .B0(cout_adj_5149), 
          .C0(n135_adj_4791), .D0(d4_adj_5676[52]), .A1(d3_adj_5675[53]), 
          .B1(cout_adj_5149), .C1(n132_adj_4790), .D1(d4_adj_5676[53]), 
          .CIN(n16310), .COUT(n16311), .S0(d4_71__N_634_adj_5692[52]), 
          .S1(d4_71__N_634_adj_5692[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_17 (.A0(d3_adj_5675[50]), .B0(cout_adj_5149), 
          .C0(n141_adj_4740), .D0(d4_adj_5676[50]), .A1(d3_adj_5675[51]), 
          .B1(cout_adj_5149), .C1(n138_adj_4741), .D1(d4_adj_5676[51]), 
          .CIN(n16309), .COUT(n16310), .S0(d4_71__N_634_adj_5692[50]), 
          .S1(d4_71__N_634_adj_5692[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_15 (.A0(d3_adj_5675[48]), .B0(cout_adj_5149), 
          .C0(n147_adj_4563), .D0(d4_adj_5676[48]), .A1(d3_adj_5675[49]), 
          .B1(cout_adj_5149), .C1(n144_adj_4739), .D1(d4_adj_5676[49]), 
          .CIN(n16308), .COUT(n16309), .S0(d4_71__N_634_adj_5692[48]), 
          .S1(d4_71__N_634_adj_5692[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_15.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[38]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[36]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    CCU2C _add_1_1493_add_4_13 (.A0(d3_adj_5675[46]), .B0(cout_adj_5149), 
          .C0(n153_adj_4561), .D0(d4_adj_5676[46]), .A1(d3_adj_5675[47]), 
          .B1(cout_adj_5149), .C1(n150_adj_4562), .D1(d4_adj_5676[47]), 
          .CIN(n16307), .COUT(n16308), .S0(d4_71__N_634_adj_5692[46]), 
          .S1(d4_71__N_634_adj_5692[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_32 (.A0(d4[30]), .B0(d3[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[31]), .B1(d3[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16070), .COUT(n16071), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_35 (.A0(d_tmp_adj_5671[68]), .B0(cout_adj_5489), 
          .C0(n87_adj_5321), .D0(n5_adj_2758), .A1(d_tmp_adj_5671[69]), 
          .B1(cout_adj_5489), .C1(n84_adj_5320), .D1(n4_adj_2759), .CIN(n16473), 
          .COUT(n16474), .S0(d6_71__N_1459_adj_5705[68]), .S1(d6_71__N_1459_adj_5705[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_29 (.A0(d7[62]), .B0(cout_adj_5050), .C0(n105_adj_4933), 
          .D0(n11_adj_4592), .A1(d7[63]), .B1(cout_adj_5050), .C1(n102_adj_4932), 
          .D1(n10_adj_4617), .CIN(n16429), .COUT(n16430), .S0(d8_71__N_1603[62]), 
          .S1(d8_71__N_1603[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_32 (.A0(d_d9_adj_5685[65]), .B0(d9_adj_5684[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[66]), .B1(d9_adj_5684[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16509), .COUT(n16510), .S0(n96_adj_4915), 
          .S1(n93_adj_4914));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_30 (.A0(d4[28]), .B0(d3[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[29]), .B1(d3[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16069), .COUT(n16070), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_30.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    CCU2C _add_1_1466_add_4_3 (.A0(d7[36]), .B0(cout_adj_5050), .C0(n183_adj_4959), 
          .D0(n37_adj_4688), .A1(d7[37]), .B1(cout_adj_5050), .C1(n180_adj_4958), 
          .D1(n36_adj_4693), .CIN(n16416), .COUT(n16417), .S0(d8_71__N_1603[36]), 
          .S1(d8_71__N_1603[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_33 (.A0(d_tmp_adj_5671[66]), .B0(cout_adj_5489), 
          .C0(n93_adj_5323), .D0(n7_adj_2756), .A1(d_tmp_adj_5671[67]), 
          .B1(cout_adj_5489), .C1(n90_adj_5322), .D1(n6_adj_2757), .CIN(n16472), 
          .COUT(n16473), .S0(d6_71__N_1459_adj_5705[66]), .S1(d6_71__N_1459_adj_5705[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_33.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    CCU2C _add_1_1481_add_4_29 (.A0(d_tmp_adj_5671[62]), .B0(cout_adj_5489), 
          .C0(n105_adj_5327), .D0(n11), .A1(d_tmp_adj_5671[63]), .B1(cout_adj_5489), 
          .C1(n102_adj_5326), .D1(n10), .CIN(n16470), .COUT(n16471), 
          .S0(d6_71__N_1459_adj_5705[62]), .S1(d6_71__N_1459_adj_5705[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_15 (.A0(d4_adj_5676[48]), .B0(cout_adj_5150), 
          .C0(n147_adj_4860), .D0(d5_adj_5677[48]), .A1(d4_adj_5676[49]), 
          .B1(cout_adj_5150), .C1(n144_adj_4859), .D1(d5_adj_5677[49]), 
          .CIN(n16352), .COUT(n16353), .S0(d5_71__N_706_adj_5693[48]), 
          .S1(d5_71__N_706_adj_5693[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_23 (.A0(d4_adj_5676[56]), .B0(cout_adj_5150), 
          .C0(n123_adj_4852), .D0(d5_adj_5677[56]), .A1(d4_adj_5676[57]), 
          .B1(cout_adj_5150), .C1(n120_adj_4851), .D1(d5_adj_5677[57]), 
          .CIN(n16356), .COUT(n16357), .S0(d5_71__N_706_adj_5693[56]), 
          .S1(d5_71__N_706_adj_5693[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_27 (.A0(d_tmp_adj_5671[60]), .B0(cout_adj_5489), 
          .C0(n111_adj_5329), .D0(n13), .A1(d_tmp_adj_5671[61]), .B1(cout_adj_5489), 
          .C1(n108_adj_5328), .D1(n12), .CIN(n16469), .COUT(n16470), 
          .S0(d6_71__N_1459_adj_5705[60]), .S1(d6_71__N_1459_adj_5705[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_25 (.A0(d_tmp_adj_5671[58]), .B0(cout_adj_5489), 
          .C0(n117_adj_5331), .D0(n15), .A1(d_tmp_adj_5671[59]), .B1(cout_adj_5489), 
          .C1(n114_adj_5330), .D1(n14), .CIN(n16468), .COUT(n16469), 
          .S0(d6_71__N_1459_adj_5705[58]), .S1(d6_71__N_1459_adj_5705[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_23 (.A0(d_tmp_adj_5671[56]), .B0(cout_adj_5489), 
          .C0(n123_adj_5333), .D0(n17), .A1(d_tmp_adj_5671[57]), .B1(cout_adj_5489), 
          .C1(n120_adj_5332), .D1(n16), .CIN(n16467), .COUT(n16468), 
          .S0(d6_71__N_1459_adj_5705[56]), .S1(d6_71__N_1459_adj_5705[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_21 (.A0(d_tmp_adj_5671[54]), .B0(cout_adj_5489), 
          .C0(n129_adj_5335), .D0(n19), .A1(d_tmp_adj_5671[55]), .B1(cout_adj_5489), 
          .C1(n126_adj_5334), .D1(n18), .CIN(n16466), .COUT(n16467), 
          .S0(d6_71__N_1459_adj_5705[54]), .S1(d6_71__N_1459_adj_5705[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_19 (.A0(d_tmp_adj_5671[52]), .B0(cout_adj_5489), 
          .C0(n135_adj_5337), .D0(n21), .A1(d_tmp_adj_5671[53]), .B1(cout_adj_5489), 
          .C1(n132_adj_5336), .D1(n20), .CIN(n16465), .COUT(n16466), 
          .S0(d6_71__N_1459_adj_5705[52]), .S1(d6_71__N_1459_adj_5705[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_19.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    CCU2C _add_1_1421_add_4_28 (.A0(d4[26]), .B0(d3[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[27]), .B1(d3[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16068), .COUT(n16069), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_26 (.A0(d4[24]), .B0(d3[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[25]), .B1(d3[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16067), .COUT(n16068), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_24 (.A0(d4[22]), .B0(d3[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[23]), .B1(d3[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16066), .COUT(n16067), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_22 (.A0(d4[20]), .B0(d3[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[21]), .B1(d3[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16065), .COUT(n16066), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_22.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i1 (.D(n126_adj_5191), .CK(CIC1_out_clkSin), .Q(ISquare[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i1.GSR = "ENABLED";
    CCU2C _add_1_1421_add_4_20 (.A0(d4[18]), .B0(d3[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[19]), .B1(d3[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16064), .COUT(n16065), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_18 (.A0(d4[16]), .B0(d3[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[17]), .B1(d3[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16063), .COUT(n16064), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_16 (.A0(d4[14]), .B0(d3[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[15]), .B1(d3[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16062), .COUT(n16063), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_14 (.A0(d4[12]), .B0(d3[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[13]), .B1(d3[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16061), .COUT(n16062), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_21 (.A0(d4_adj_5676[54]), .B0(cout_adj_5150), 
          .C0(n129_adj_4854), .D0(d5_adj_5677[54]), .A1(d4_adj_5676[55]), 
          .B1(cout_adj_5150), .C1(n126_adj_4853), .D1(d5_adj_5677[55]), 
          .CIN(n16355), .COUT(n16356), .S0(d5_71__N_706_adj_5693[54]), 
          .S1(d5_71__N_706_adj_5693[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_12 (.A0(d4[10]), .B0(d3[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[11]), .B1(d3[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16060), .COUT(n16061), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_10 (.A0(d4[8]), .B0(d3[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[9]), .B1(d3[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16059), .COUT(n16060), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_8 (.A0(d4[6]), .B0(d3[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[7]), .B1(d3[7]), .C1(GND_net), .D1(VCC_net), .CIN(n16058), 
          .COUT(n16059), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_6 (.A0(d4[4]), .B0(d3[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[5]), .B1(d3[5]), .C1(GND_net), .D1(VCC_net), .CIN(n16057), 
          .COUT(n16058), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_6 (.A0(d4_adj_5676[39]), .B0(d3_adj_5675[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[40]), .B1(d3_adj_5675[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16269), .COUT(n16270), .S0(n174_adj_4554), 
          .S1(n171_adj_4555));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_4 (.A0(d4_adj_5676[37]), .B0(d3_adj_5675[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[38]), .B1(d3_adj_5675[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16268), .COUT(n16269), .S0(n180_adj_4552), 
          .S1(n177_adj_4553));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_26 (.A0(d4_adj_5676[59]), .B0(d3_adj_5675[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[60]), .B1(d3_adj_5675[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16279), .COUT(n16280), .S0(n114_adj_4744), 
          .S1(n111_adj_4742));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_26.INJECT1_1 = "NO";
    LUT4 i2342_3_lut_4_lut (.A(n18267), .B(n18138), .C(n18268), .D(n136), 
         .Z(n12057)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2342_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_326_i25_4_lut (.A(n11995), .B(n247_adj_5429), .C(n18135), 
         .D(n2593), .Z(n2368)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i25_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1490_add_4_19 (.A0(d4_adj_5676[52]), .B0(cout_adj_5150), 
          .C0(n135_adj_4856), .D0(d5_adj_5677[52]), .A1(d4_adj_5676[53]), 
          .B1(cout_adj_5150), .C1(n132_adj_4855), .D1(d5_adj_5677[53]), 
          .CIN(n16354), .COUT(n16355), .S0(d5_71__N_706_adj_5693[52]), 
          .S1(d5_71__N_706_adj_5693[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_35 (.A0(d7[68]), .B0(cout_adj_5050), .C0(n87_adj_4927), 
          .D0(n5_adj_4689), .A1(d7[69]), .B1(cout_adj_5050), .C1(n84_adj_4926), 
          .D1(n4_adj_4690), .CIN(n16432), .COUT(n16433), .S0(d8_71__N_1603[68]), 
          .S1(d8_71__N_1603[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5050), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16416));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1466_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1466_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_1.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i0 (.D(n321), .CK(clk_80mhz), .Q(phase_accum_adj_5665[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1421_add_4_4 (.A0(d4[2]), .B0(d3[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[3]), .B1(d3[3]), .C1(GND_net), .D1(VCC_net), .CIN(n16056), 
          .COUT(n16057), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_4.INJECT1_1 = "NO";
    LUT4 mux_326_i26_4_lut (.A(n8_adj_5661), .B(n244_adj_5428), .C(n18135), 
         .D(n17322), .Z(n2367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i26_4_lut.init = 16'hcfca;
    LUT4 i2334_3_lut_4_lut (.A(n18267), .B(n18138), .C(led_c_3), .D(n151), 
         .Z(n12049)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2334_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1484_add_4_37 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16412), .S0(n76));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1484_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_11 (.A0(d3_adj_5675[44]), .B0(cout_adj_5149), 
          .C0(n159_adj_4559), .D0(d4_adj_5676[44]), .A1(d3_adj_5675[45]), 
          .B1(cout_adj_5149), .C1(n156_adj_4560), .D1(d4_adj_5676[45]), 
          .CIN(n16306), .COUT(n16307), .S0(d4_71__N_634_adj_5692[44]), 
          .S1(d4_71__N_634_adj_5692[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_13 (.A0(d4_adj_5676[46]), .B0(cout_adj_5150), 
          .C0(n153_adj_4862), .D0(d5_adj_5677[46]), .A1(d4_adj_5676[47]), 
          .B1(cout_adj_5150), .C1(n150_adj_4861), .D1(d5_adj_5677[47]), 
          .CIN(n16351), .COUT(n16352), .S0(d5_71__N_706_adj_5693[46]), 
          .S1(d5_71__N_706_adj_5693[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_13.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_159_4_lut (.A(led_c_4), .B(n18145), .C(n18144), 
         .D(n26_adj_5659), .Z(n18129)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_rep_159_4_lut.init = 16'hf400;
    CCU2C _add_1_1421_add_4_2 (.A0(d4[0]), .B0(d3[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[1]), .B1(d3[1]), .C1(GND_net), .D1(VCC_net), .COUT(n16056), 
          .S1(d4_71__N_634[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1421_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_27 (.A0(d7[60]), .B0(cout_adj_5050), .C0(n111_adj_4935), 
          .D0(n13_adj_4576), .A1(d7[61]), .B1(cout_adj_5050), .C1(n108_adj_4934), 
          .D1(n12_adj_4577), .CIN(n16428), .COUT(n16429), .S0(d8_71__N_1603[60]), 
          .S1(d8_71__N_1603[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_25 (.A0(d7[58]), .B0(cout_adj_5050), .C0(n117_adj_4937), 
          .D0(n15_adj_4573), .A1(d7[59]), .B1(cout_adj_5050), .C1(n114_adj_4936), 
          .D1(n14_adj_4575), .CIN(n16427), .COUT(n16428), .S0(d8_71__N_1603[58]), 
          .S1(d8_71__N_1603[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_23 (.A0(d7[56]), .B0(cout_adj_5050), .C0(n123_adj_4939), 
          .D0(n17_adj_4571), .A1(d7[57]), .B1(cout_adj_5050), .C1(n120_adj_4938), 
          .D1(n16_adj_4572), .CIN(n16426), .COUT(n16427), .S0(d8_71__N_1603[56]), 
          .S1(d8_71__N_1603[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_28 (.A0(d4_adj_5676[26]), .B0(d3_adj_5675[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[27]), .B1(d3_adj_5675[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16489), .COUT(n16490), .S0(d4_71__N_634_adj_5692[26]), 
          .S1(d4_71__N_634_adj_5692[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4_adj_5676[36]), .B1(d3_adj_5675[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16268), .S1(n183_adj_4551));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1577_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_26 (.A0(d4_adj_5676[24]), .B0(d3_adj_5675[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[25]), .B1(d3_adj_5675[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16488), .COUT(n16489), .S0(d4_71__N_634_adj_5692[24]), 
          .S1(d4_71__N_634_adj_5692[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_26.INJECT1_1 = "NO";
    LUT4 i6624_4_lut (.A(n26_adj_5659), .B(n18267), .C(n18191), .D(n18144), 
         .Z(n13099)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i6624_4_lut.init = 16'h575f;
    LUT4 led_c_4_bdd_4_lut (.A(led_c_2), .B(led_c_0), .C(led_c_1), .D(n18268), 
         .Z(n18086)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B+(C (D)+!C !(D)))) */ ;
    defparam led_c_4_bdd_4_lut.init = 16'ha9b0;
    LUT4 n18086_bdd_2_lut (.A(n18086), .B(led_c_4), .Z(n18087)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n18086_bdd_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_57 (.A(led_c_4), .B(n18142), .C(led_c_3), 
         .D(led_c_2), .Z(n17310)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_57.init = 16'hfeff;
    LUT4 i6642_4_lut_rep_217 (.A(n17593), .B(n18142), .C(n18087), .D(n17963), 
         .Z(n18301)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i6642_4_lut_rep_217.init = 16'h3032;
    CCU2C _add_1_1586_add_4_38 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16267), .S0(n78_adj_5035));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1586_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_38.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(led_c_3), .B(n238), .Z(n8_adj_5661)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i6642_4_lut_rep_218 (.A(n17593), .B(n18142), .C(n18087), .D(n17963), 
         .Z(clk_80mhz_enable_881)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i6642_4_lut_rep_218.init = 16'h3032;
    CCU2C _add_1_1481_add_4_17 (.A0(d_tmp_adj_5671[50]), .B0(cout_adj_5489), 
          .C0(n141_adj_5339), .D0(n23_adj_2755), .A1(d_tmp_adj_5671[51]), 
          .B1(cout_adj_5489), .C1(n138_adj_5338), .D1(n22), .CIN(n16464), 
          .COUT(n16465), .S0(d6_71__N_1459_adj_5705[50]), .S1(d6_71__N_1459_adj_5705[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_37 (.A0(d_tmp[70]), .B0(cout_adj_5496), .C0(n81_adj_5052), 
          .D0(n3_adj_4767), .A1(d_tmp[71]), .B1(cout_adj_5496), .C1(n78_adj_5051), 
          .D1(n2_adj_4768), .CIN(n16341), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_24 (.A0(d4_adj_5676[22]), .B0(d3_adj_5675[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[23]), .B1(d3_adj_5675[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16487), .COUT(n16488), .S0(d4_71__N_634_adj_5692[22]), 
          .S1(d4_71__N_634_adj_5692[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_24.INJECT1_1 = "NO";
    LUT4 n17536_bdd_4_lut (.A(n17536), .B(n17298), .C(n18267), .D(n26_adj_5659), 
         .Z(n2845)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n17536_bdd_4_lut.init = 16'hca00;
    CCU2C _add_1_1481_add_4_13 (.A0(d_tmp_adj_5671[46]), .B0(cout_adj_5489), 
          .C0(n153_adj_5343), .D0(n27_adj_2751), .A1(d_tmp_adj_5671[47]), 
          .B1(cout_adj_5489), .C1(n150_adj_5342), .D1(n26_adj_2752), .CIN(n16462), 
          .COUT(n16463), .S0(d6_71__N_1459_adj_5705[46]), .S1(d6_71__N_1459_adj_5705[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_14 (.A0(d_d9_adj_5685[47]), .B0(d9_adj_5684[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[48]), .B1(d9_adj_5684[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16500), .COUT(n16501));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_3 (.A0(d4_adj_5676[36]), .B0(cout_adj_5150), 
          .C0(n183_adj_4872), .D0(d5_adj_5677[36]), .A1(d4_adj_5676[37]), 
          .B1(cout_adj_5150), .C1(n180_adj_4871), .D1(d5_adj_5677[37]), 
          .CIN(n16346), .COUT(n16347), .S0(d5_71__N_706_adj_5693[36]), 
          .S1(d5_71__N_706_adj_5693[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_12 (.A0(d_d9_adj_5685[45]), .B0(d9_adj_5684[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[46]), .B1(d9_adj_5684[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16499), .COUT(n16500));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_36 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16266), .COUT(n16267), .S0(n84_adj_5037), .S1(n81_adj_5036));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_36.INJECT1_1 = "NO";
    FD1S3AX _add_1_1649_i7 (.D(cout_adj_4997), .CK(clk_80mhz), .Q(PWMOutP4_c));
    defparam _add_1_1649_i7.GSR = "ENABLED";
    OB led_pad_6 (.I(led_c_6), .O(led[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    CCU2C _add_1_1496_add_4_37 (.A0(d2_adj_5674[70]), .B0(cout_adj_5132), 
          .C0(n81_adj_5624), .D0(d3_adj_5675[70]), .A1(d2_adj_5674[71]), 
          .B1(cout_adj_5132), .C1(n78_adj_5623), .D1(d3_adj_5675[71]), 
          .CIN(n16053), .S0(d3_71__N_562_adj_5691[70]), .S1(d3_71__N_562_adj_5691[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_34 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16265), .COUT(n16266), .S0(n90_adj_5039), .S1(n87_adj_5038));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_32 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16264), .COUT(n16265), .S0(n96_adj_5041), .S1(n93_adj_5040));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_30 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16263), .COUT(n16264), .S0(n102_adj_5043), .S1(n99_adj_5042));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_28 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16262), .COUT(n16263), .S0(n108_adj_5045), .S1(n105_adj_5044));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_26 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16261), .COUT(n16262), .S0(n114_adj_5047), .S1(n111_adj_5046));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_24 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16260), .COUT(n16261), .S0(n120_adj_5049), .S1(n117_adj_5048));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_7 (.A0(d4_adj_5676[40]), .B0(cout_adj_5150), 
          .C0(n171_adj_4868), .D0(d5_adj_5677[40]), .A1(d4_adj_5676[41]), 
          .B1(cout_adj_5150), .C1(n168_adj_4867), .D1(d5_adj_5677[41]), 
          .CIN(n16348), .COUT(n16349), .S0(d5_71__N_706_adj_5693[40]), 
          .S1(d5_71__N_706_adj_5693[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_7.INJECT1_1 = "NO";
    OB led_pad_7 (.I(led_c_7), .O(led[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    CCU2C _add_1_1586_add_4_22 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16259), .COUT(n16260));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_20 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16258), .COUT(n16259));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_18 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16257), .COUT(n16258));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_16 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16256), .COUT(n16257));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_14 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16255), .COUT(n16256));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_22 (.A0(d4_adj_5676[20]), .B0(d3_adj_5675[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[21]), .B1(d3_adj_5675[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16486), .COUT(n16487), .S0(d4_71__N_634_adj_5692[20]), 
          .S1(d4_71__N_634_adj_5692[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_12 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16254), .COUT(n16255));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_10 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16253), .COUT(n16254));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_36 (.A0(d4_adj_5676[69]), .B0(d3_adj_5675[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[70]), .B1(d3_adj_5675[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16284), .COUT(n16285), .S0(n84), 
          .S1(n81));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_8 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16252), .COUT(n16253));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_20 (.A0(d4_adj_5676[18]), .B0(d3_adj_5675[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[19]), .B1(d3_adj_5675[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16485), .COUT(n16486), .S0(d4_71__N_634_adj_5692[18]), 
          .S1(d4_71__N_634_adj_5692[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_35 (.A0(d_tmp[68]), .B0(cout_adj_5496), .C0(n87_adj_5054), 
          .D0(n5_adj_4765), .A1(d_tmp[69]), .B1(cout_adj_5496), .C1(n84_adj_5053), 
          .D1(n4_adj_4766), .CIN(n16340), .COUT(n16341), .S0(d6_71__N_1459[68]), 
          .S1(d6_71__N_1459[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_6 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16251), .COUT(n16252));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_4 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16250), .COUT(n16251));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16250));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1586_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1586_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_20 (.A0(n912), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16249), .S0(d_out_d_11__N_2335[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_20.INIT0 = 16'h555f;
    defparam _add_1_1589_add_4_20.INIT1 = 16'h0000;
    defparam _add_1_1589_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_20.INJECT1_1 = "NO";
    LUT4 i349_2_lut_rep_165_4_lut (.A(n26_adj_5659), .B(n18145), .C(led_c_4), 
         .D(n18268), .Z(n18135)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i349_2_lut_rep_165_4_lut.init = 16'h0080;
    CCU2C _add_1_1589_add_4_18 (.A0(ISquare[31]), .B0(n914), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n913), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16248), .COUT(n16249));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_11 (.A0(d4_adj_5676[44]), .B0(cout_adj_5150), 
          .C0(n159_adj_4864), .D0(d5_adj_5677[44]), .A1(d4_adj_5676[45]), 
          .B1(cout_adj_5150), .C1(n156_adj_4863), .D1(d5_adj_5677[45]), 
          .CIN(n16350), .COUT(n16351), .S0(d5_71__N_706_adj_5693[44]), 
          .S1(d5_71__N_706_adj_5693[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_10 (.A0(d_d9_adj_5685[43]), .B0(d9_adj_5684[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[44]), .B1(d9_adj_5684[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16498), .COUT(n16499));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_33 (.A0(d_tmp[66]), .B0(cout_adj_5496), .C0(n93_adj_5056), 
          .D0(n7_adj_4763), .A1(d_tmp[67]), .B1(cout_adj_5496), .C1(n90_adj_5055), 
          .D1(n6_adj_4764), .CIN(n16339), .COUT(n16340), .S0(d6_71__N_1459[66]), 
          .S1(d6_71__N_1459[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_16 (.A0(n916), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n915), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16247), .COUT(n16248));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1589_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_14 (.A0(d_out_d_11__N_1874[17]), .B0(n918), 
          .C0(GND_net), .D0(VCC_net), .A1(ISquare[31]), .B1(n18150), 
          .C1(n917), .D1(VCC_net), .CIN(n16246), .COUT(n16247));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_1589_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_12 (.A0(d_out_d_11__N_1878[17]), .B0(n920), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n919), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16245), .COUT(n16246));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_12.INJECT1_1 = "NO";
    OB o_Tx_Serial_pad (.I(GND_net), .O(o_Tx_Serial));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(48[11:22])
    CCU2C _add_1_1589_add_4_10 (.A0(d_out_d_11__N_1882[17]), .B0(n922), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n921), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16244), .COUT(n16245));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_10.INJECT1_1 = "NO";
    \uart_rx(CLKS_PER_BIT=87)  uart_rx1 (.clk_80mhz(clk_80mhz), .i_Rx_Serial_c(i_Rx_Serial_c), 
            .o_Rx_Byte1({o_Rx_Byte1}), .GND_net(GND_net), .VCC_net(VCC_net), 
            .o_Rx_DV1(o_Rx_DV1)) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(230[32] 235[2])
    CCU2C _add_1_1589_add_4_8 (.A0(d_out_d_11__N_1886[17]), .B0(n924), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n923), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16243), .COUT(n16244));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_8.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_169_3_lut (.A(led_c_6), .B(n18149), .C(led_c_4), 
         .Z(n18139)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_2_lut_rep_169_3_lut.init = 16'hfdfd;
    CCU2C _add_1_1589_add_4_6 (.A0(d_out_d_11__N_1890[17]), .B0(n926), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n925), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16242), .COUT(n16243));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_6.INJECT1_1 = "NO";
    OB led_pad_5 (.I(led_c_5), .O(led[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    CCU2C _add_1_1493_add_4_9 (.A0(d3_adj_5675[42]), .B0(cout_adj_5149), 
          .C0(n165_adj_4557), .D0(d4_adj_5676[42]), .A1(d3_adj_5675[43]), 
          .B1(cout_adj_5149), .C1(n162_adj_4558), .D1(d4_adj_5676[43]), 
          .CIN(n16305), .COUT(n16306), .S0(d4_71__N_634_adj_5692[42]), 
          .S1(d4_71__N_634_adj_5692[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_9.INJECT1_1 = "NO";
    LUT4 i26_4_lut (.A(n2593), .B(n253_adj_5431), .C(n18135), .D(n13_adj_5485), 
         .Z(n11_adj_5484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i26_4_lut.init = 16'hcacf;
    CCU2C _add_1_1484_add_4_35 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16411), .COUT(n16412), .S0(n82), .S1(n79));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_35.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i8 (.D(o_Rx_Byte1[7]), .CK(clk_80mhz), .Q(led_c_7));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i8.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i7 (.D(o_Rx_Byte1[6]), .CK(clk_80mhz), .Q(led_c_6));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i6 (.D(o_Rx_Byte1[5]), .CK(clk_80mhz), .Q(led_c_5));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i5 (.D(o_Rx_Byte1[4]), .CK(clk_80mhz), .Q(led_c_4));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i4 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(led_c_3));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i3 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(led_c_2));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i2 (.D(o_Rx_Byte1[1]), .CK(clk_80mhz), .Q(led_c_1));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    CCU2C _add_1_1493_add_4_7 (.A0(d3_adj_5675[40]), .B0(cout_adj_5149), 
          .C0(n171_adj_4555), .D0(d4_adj_5676[40]), .A1(d3_adj_5675[41]), 
          .B1(cout_adj_5149), .C1(n168_adj_4556), .D1(d4_adj_5676[41]), 
          .CIN(n16304), .COUT(n16305), .S0(d4_71__N_634_adj_5692[40]), 
          .S1(d4_71__N_634_adj_5692[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_4 (.A0(d_out_d_11__N_1892[17]), .B0(ISquare[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1892[17]), .B1(n927), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16241), .COUT(n16242));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_5 (.A0(d3_adj_5675[38]), .B0(cout_adj_5149), 
          .C0(n177_adj_4553), .D0(d4_adj_5676[38]), .A1(d3_adj_5675[39]), 
          .B1(cout_adj_5149), .C1(n174_adj_4554), .D1(d4_adj_5676[39]), 
          .CIN(n16303), .COUT(n16304), .S0(d4_71__N_634_adj_5692[38]), 
          .S1(d4_71__N_634_adj_5692[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_3 (.A0(d3_adj_5675[36]), .B0(cout_adj_5149), 
          .C0(n183_adj_4551), .D0(d4_adj_5676[36]), .A1(d3_adj_5675[37]), 
          .B1(cout_adj_5149), .C1(n180_adj_4552), .D1(d4_adj_5676[37]), 
          .CIN(n16302), .COUT(n16303), .S0(d4_71__N_634_adj_5692[36]), 
          .S1(d4_71__N_634_adj_5692[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5149), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16302));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1493_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1493_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_1.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_26 (.A0(MultResult2[23]), .B0(MultResult1[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16298), .S0(n54_adj_5167));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_26.INIT0 = 16'h666a;
    defparam ISquare_add_4_26.INIT1 = 16'h0000;
    defparam ISquare_add_4_26.INJECT1_0 = "NO";
    defparam ISquare_add_4_26.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_24 (.A0(MultResult2[22]), .B0(MultResult1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[23]), .B1(MultResult1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16297), .COUT(n16298), .S0(n60_adj_5169), 
          .S1(n57_adj_5168));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_24.INIT0 = 16'h666a;
    defparam ISquare_add_4_24.INIT1 = 16'h666a;
    defparam ISquare_add_4_24.INJECT1_0 = "NO";
    defparam ISquare_add_4_24.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_22 (.A0(MultResult2[20]), .B0(MultResult1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[21]), .B1(MultResult1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16296), .COUT(n16297), .S0(n66_adj_5171), 
          .S1(n63_adj_5170));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_22.INIT0 = 16'h666a;
    defparam ISquare_add_4_22.INIT1 = 16'h666a;
    defparam ISquare_add_4_22.INJECT1_0 = "NO";
    defparam ISquare_add_4_22.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_20 (.A0(MultResult2[18]), .B0(MultResult1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[19]), .B1(MultResult1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16295), .COUT(n16296), .S0(n72_adj_5173), 
          .S1(n69_adj_5172));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_20.INIT0 = 16'h666a;
    defparam ISquare_add_4_20.INIT1 = 16'h666a;
    defparam ISquare_add_4_20.INJECT1_0 = "NO";
    defparam ISquare_add_4_20.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_18 (.A0(MultResult2[16]), .B0(MultResult1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[17]), .B1(MultResult1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16294), .COUT(n16295), .S0(n78_adj_5175), 
          .S1(n75_adj_5174));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_18.INIT0 = 16'h666a;
    defparam ISquare_add_4_18.INIT1 = 16'h666a;
    defparam ISquare_add_4_18.INJECT1_0 = "NO";
    defparam ISquare_add_4_18.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_16 (.A0(MultResult2[14]), .B0(MultResult1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[15]), .B1(MultResult1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16293), .COUT(n16294), .S0(n84_adj_5177), 
          .S1(n81_adj_5176));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_16.INIT0 = 16'h666a;
    defparam ISquare_add_4_16.INIT1 = 16'h666a;
    defparam ISquare_add_4_16.INJECT1_0 = "NO";
    defparam ISquare_add_4_16.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_14 (.A0(MultResult2[12]), .B0(MultResult1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[13]), .B1(MultResult1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16292), .COUT(n16293), .S0(n90_adj_5179), 
          .S1(n87_adj_5178));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_14.INIT0 = 16'h666a;
    defparam ISquare_add_4_14.INIT1 = 16'h666a;
    defparam ISquare_add_4_14.INJECT1_0 = "NO";
    defparam ISquare_add_4_14.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_12 (.A0(MultResult2[10]), .B0(MultResult1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[11]), .B1(MultResult1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16291), .COUT(n16292), .S0(n96_adj_5181), 
          .S1(n93_adj_5180));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_12.INIT0 = 16'h666a;
    defparam ISquare_add_4_12.INIT1 = 16'h666a;
    defparam ISquare_add_4_12.INJECT1_0 = "NO";
    defparam ISquare_add_4_12.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_10 (.A0(MultResult2[8]), .B0(MultResult1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[9]), .B1(MultResult1[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16290), .COUT(n16291), .S0(n102_adj_5183), 
          .S1(n99_adj_5182));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_10.INIT0 = 16'h666a;
    defparam ISquare_add_4_10.INIT1 = 16'h666a;
    defparam ISquare_add_4_10.INJECT1_0 = "NO";
    defparam ISquare_add_4_10.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_8 (.A0(MultResult2[6]), .B0(MultResult1[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[7]), .B1(MultResult1[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16289), .COUT(n16290), .S0(n108_adj_5185), 
          .S1(n105_adj_5184));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_8.INIT0 = 16'h666a;
    defparam ISquare_add_4_8.INIT1 = 16'h666a;
    defparam ISquare_add_4_8.INJECT1_0 = "NO";
    defparam ISquare_add_4_8.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_6 (.A0(MultResult2[4]), .B0(MultResult1[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[5]), .B1(MultResult1[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16288), .COUT(n16289), .S0(n114_adj_5187), 
          .S1(n111_adj_5186));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_6.INIT0 = 16'h666a;
    defparam ISquare_add_4_6.INIT1 = 16'h666a;
    defparam ISquare_add_4_6.INJECT1_0 = "NO";
    defparam ISquare_add_4_6.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_4 (.A0(MultResult2[2]), .B0(MultResult1[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[3]), .B1(MultResult1[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16287), .COUT(n16288), .S0(n120_adj_5189), 
          .S1(n117_adj_5188));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_4.INIT0 = 16'h666a;
    defparam ISquare_add_4_4.INIT1 = 16'h666a;
    defparam ISquare_add_4_4.INJECT1_0 = "NO";
    defparam ISquare_add_4_4.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_2 (.A0(MultResult2[0]), .B0(MultResult1[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[1]), .B1(MultResult1[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16287), .S1(n123_adj_5190));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_2.INIT0 = 16'h0008;
    defparam ISquare_add_4_2.INIT1 = 16'h666a;
    defparam ISquare_add_4_2.INJECT1_0 = "NO";
    defparam ISquare_add_4_2.INJECT1_1 = "NO";
    LUT4 i2320_3_lut_4_lut (.A(n18138), .B(n18267), .C(n18268), .D(n175), 
         .Z(n12035)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2320_3_lut_4_lut.init = 16'hf707;
    CCU2C _add_1_1577_add_4_38 (.A0(d4_adj_5676[71]), .B0(d3_adj_5675[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16285), .S0(n78));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1577_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16241));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1589_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1589_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_2.INJECT1_1 = "NO";
    LUT4 mux_326_i24_4_lut (.A(n11993), .B(n250_adj_5430), .C(n18135), 
         .D(n2593), .Z(n2369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i24_4_lut.init = 16'hcfca;
    LUT4 i1_4_lut (.A(led_c_5), .B(led_c_7), .C(led_c_6), .D(o_Rx_DV), 
         .Z(n26_adj_5659)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_4_lut.init = 16'h2000;
    FD1P3AX phase_inc_carrGen_i0_i1 (.D(n320), .SP(clk_80mhz_enable_831), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    OB led_pad_4 (.I(led_c_4), .O(led[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    OB led_pad_3 (.I(led_c_3), .O(led[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    OB led_pad_2 (.I(led_c_2), .O(led[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    OB led_pad_1 (.I(led_c_1), .O(led[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    OB led_pad_0 (.I(led_c_0), .O(led[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(49[18:21])
    OB XOut_pad (.I(GND_net), .O(XOut));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(53[9:13])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(55[9:16])
    OB PWMOut_pad (.I(PWMOutP4_c), .O(PWMOut));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(56[9:15])
    OB PWMOutP1_pad (.I(PWMOutP4_c), .O(PWMOutP1));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(57[9:17])
    OB PWMOutP2_pad (.I(PWMOutP4_c), .O(PWMOutP2));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(58[9:17])
    OB PWMOutP3_pad (.I(PWMOutP4_c), .O(PWMOutP3));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(59[9:17])
    OB PWMOutP4_pad (.I(PWMOutP4_c), .O(PWMOutP4));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(60[9:17])
    OB PWMOutN1_pad (.I(PWMOutN4_c), .O(PWMOutN1));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(61[9:17])
    OB PWMOutN2_pad (.I(PWMOutN4_c), .O(PWMOutN2));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(62[9:17])
    OB PWMOutN3_pad (.I(PWMOutN4_c), .O(PWMOutN3));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(63[9:17])
    OB PWMOutN4_pad (.I(PWMOutN4_c), .O(PWMOutN4));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(64[9:17])
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(65[9:15])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(66[9:16])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(67[9:23])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(47[13:24])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(54[9:13])
    IB clk_25mhz_pad (.I(clk_25mhz), .O(clk_25mhz_c));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(68[8:17])
    CCU2C _add_1_1484_add_4_33 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16410), .COUT(n16411), .S0(n88), .S1(n85));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_31 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16409), .COUT(n16410), .S0(n94), .S1(n91));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_29 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16408), .COUT(n16409), .S0(n100), .S1(n97));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_27 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16407), .COUT(n16408), .S0(n106), .S1(n103));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_25 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16406), .COUT(n16407), .S0(n112), .S1(n109));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_23 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16405), .COUT(n16406), .S0(n118), .S1(n115));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_21 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16404), .COUT(n16405));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_19 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16403), .COUT(n16404));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_17 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16402), .COUT(n16403));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_15 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16401), .COUT(n16402));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_13 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16400), .COUT(n16401));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_11 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16399), .COUT(n16400));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_9 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16398), .COUT(n16399));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_7 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16397), .COUT(n16398));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_5 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16396), .COUT(n16397));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_3 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16395), .COUT(n16396));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16395));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1484_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_17 (.A0(count_adj_5688[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16394), .S0(n36_adj_5151));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1445_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_15 (.A0(count_adj_5688[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16393), .COUT(n16394), .S0(n42_adj_5153), 
          .S1(n39_adj_5152));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_13 (.A0(count_adj_5688[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16392), .COUT(n16393), .S0(n48_adj_5155), 
          .S1(n45_adj_5154));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_11 (.A0(count_adj_5688[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16391), .COUT(n16392), .S0(n54_adj_5157), 
          .S1(n51_adj_5156));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_9 (.A0(count_adj_5688[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16390), .COUT(n16391), .S0(n60_adj_5159), 
          .S1(n57_adj_5158));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_7 (.A0(count_adj_5688[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16389), .COUT(n16390), .S0(n66_adj_5161), 
          .S1(n63_adj_5160));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_5 (.A0(count_adj_5688[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16388), .COUT(n16389), .S0(n72_adj_5163), 
          .S1(n69_adj_5162));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_3 (.A0(count_adj_5688[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5688[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16387), .COUT(n16388), .S0(n78_adj_5165), 
          .S1(n75_adj_5164));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_adj_5688[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16387), .S1(n81_adj_5166));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1445_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1445_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_37 (.A0(d8[70]), .B0(cout_adj_4998), .C0(n81_adj_5000), 
          .D0(n3_adj_4834), .A1(d8[71]), .B1(cout_adj_4998), .C1(n78_adj_4999), 
          .D1(n2_adj_4835), .CIN(n16385), .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_35 (.A0(d8[68]), .B0(cout_adj_4998), .C0(n87_adj_5002), 
          .D0(n5_adj_4832), .A1(d8[69]), .B1(cout_adj_4998), .C1(n84_adj_5001), 
          .D1(n4_adj_4833), .CIN(n16384), .COUT(n16385), .S0(d9_71__N_1675[68]), 
          .S1(d9_71__N_1675[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_33 (.A0(d8[66]), .B0(cout_adj_4998), .C0(n93_adj_5004), 
          .D0(n7_adj_4830), .A1(d8[67]), .B1(cout_adj_4998), .C1(n90_adj_5003), 
          .D1(n6_adj_4831), .CIN(n16383), .COUT(n16384), .S0(d9_71__N_1675[66]), 
          .S1(d9_71__N_1675[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_31 (.A0(d8[64]), .B0(cout_adj_4998), .C0(n99_adj_5006), 
          .D0(n9_adj_4828), .A1(d8[65]), .B1(cout_adj_4998), .C1(n96_adj_5005), 
          .D1(n8_adj_4829), .CIN(n16382), .COUT(n16383), .S0(d9_71__N_1675[64]), 
          .S1(d9_71__N_1675[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_29 (.A0(d8[62]), .B0(cout_adj_4998), .C0(n105_adj_5008), 
          .D0(n11_adj_4826), .A1(d8[63]), .B1(cout_adj_4998), .C1(n102_adj_5007), 
          .D1(n10_adj_4827), .CIN(n16381), .COUT(n16382), .S0(d9_71__N_1675[62]), 
          .S1(d9_71__N_1675[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_27 (.A0(d8[60]), .B0(cout_adj_4998), .C0(n111_adj_5010), 
          .D0(n13_adj_4824), .A1(d8[61]), .B1(cout_adj_4998), .C1(n108_adj_5009), 
          .D1(n12_adj_4825), .CIN(n16380), .COUT(n16381), .S0(d9_71__N_1675[60]), 
          .S1(d9_71__N_1675[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_25 (.A0(d8[58]), .B0(cout_adj_4998), .C0(n117_adj_5012), 
          .D0(n15_adj_4822), .A1(d8[59]), .B1(cout_adj_4998), .C1(n114_adj_5011), 
          .D1(n14_adj_4823), .CIN(n16379), .COUT(n16380), .S0(d9_71__N_1675[58]), 
          .S1(d9_71__N_1675[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_23 (.A0(d8[56]), .B0(cout_adj_4998), .C0(n123_adj_5014), 
          .D0(n17_adj_4820), .A1(d8[57]), .B1(cout_adj_4998), .C1(n120_adj_5013), 
          .D1(n16_adj_4821), .CIN(n16378), .COUT(n16379), .S0(d9_71__N_1675[56]), 
          .S1(d9_71__N_1675[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_21 (.A0(d8[54]), .B0(cout_adj_4998), .C0(n129_adj_5016), 
          .D0(n19_adj_4818), .A1(d8[55]), .B1(cout_adj_4998), .C1(n126_adj_5015), 
          .D1(n18_adj_4819), .CIN(n16377), .COUT(n16378), .S0(d9_71__N_1675[54]), 
          .S1(d9_71__N_1675[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_19 (.A0(d8[52]), .B0(cout_adj_4998), .C0(n135_adj_5018), 
          .D0(n21_adj_4816), .A1(d8[53]), .B1(cout_adj_4998), .C1(n132_adj_5017), 
          .D1(n20_adj_4817), .CIN(n16376), .COUT(n16377), .S0(d9_71__N_1675[52]), 
          .S1(d9_71__N_1675[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_17 (.A0(d8[50]), .B0(cout_adj_4998), .C0(n141_adj_5020), 
          .D0(n23_adj_4814), .A1(d8[51]), .B1(cout_adj_4998), .C1(n138_adj_5019), 
          .D1(n22_adj_4815), .CIN(n16375), .COUT(n16376), .S0(d9_71__N_1675[50]), 
          .S1(d9_71__N_1675[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_15 (.A0(d8[48]), .B0(cout_adj_4998), .C0(n147_adj_5022), 
          .D0(n25_adj_4782), .A1(d8[49]), .B1(cout_adj_4998), .C1(n144_adj_5021), 
          .D1(n24_adj_4783), .CIN(n16374), .COUT(n16375), .S0(d9_71__N_1675[48]), 
          .S1(d9_71__N_1675[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_13 (.A0(d8[46]), .B0(cout_adj_4998), .C0(n153_adj_5024), 
          .D0(n27_adj_4780), .A1(d8[47]), .B1(cout_adj_4998), .C1(n150_adj_5023), 
          .D1(n26_adj_4781), .CIN(n16373), .COUT(n16374), .S0(d9_71__N_1675[46]), 
          .S1(d9_71__N_1675[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_11 (.A0(d8[44]), .B0(cout_adj_4998), .C0(n159_adj_5026), 
          .D0(n29_adj_4778), .A1(d8[45]), .B1(cout_adj_4998), .C1(n156_adj_5025), 
          .D1(n28_adj_4779), .CIN(n16372), .COUT(n16373), .S0(d9_71__N_1675[44]), 
          .S1(d9_71__N_1675[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_9 (.A0(d8[42]), .B0(cout_adj_4998), .C0(n165_adj_5028), 
          .D0(n31_adj_4776), .A1(d8[43]), .B1(cout_adj_4998), .C1(n162_adj_5027), 
          .D1(n30_adj_4777), .CIN(n16371), .COUT(n16372), .S0(d9_71__N_1675[42]), 
          .S1(d9_71__N_1675[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_7 (.A0(d8[40]), .B0(cout_adj_4998), .C0(n171_adj_5030), 
          .D0(n33_adj_4774), .A1(d8[41]), .B1(cout_adj_4998), .C1(n168_adj_5029), 
          .D1(n32_adj_4775), .CIN(n16370), .COUT(n16371), .S0(d9_71__N_1675[40]), 
          .S1(d9_71__N_1675[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_5 (.A0(d8[38]), .B0(cout_adj_4998), .C0(n177_adj_5032), 
          .D0(n35_adj_4772), .A1(d8[39]), .B1(cout_adj_4998), .C1(n174_adj_5031), 
          .D1(n34_adj_4773), .CIN(n16369), .COUT(n16370), .S0(d9_71__N_1675[38]), 
          .S1(d9_71__N_1675[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_3 (.A0(d8[36]), .B0(cout_adj_4998), .C0(n183_adj_5034), 
          .D0(n37_adj_4770), .A1(d8[37]), .B1(cout_adj_4998), .C1(n180_adj_5033), 
          .D1(n36_adj_4771), .CIN(n16368), .COUT(n16369), .S0(d9_71__N_1675[36]), 
          .S1(d9_71__N_1675[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_8 (.A0(d_d9_adj_5685[41]), .B0(d9_adj_5684[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[42]), .B1(d9_adj_5684[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16497), .COUT(n16498));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_8.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[56]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[58]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[60]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[62]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    LUT4 i1_4_lut_then_3_lut (.A(led_c_3), .B(led_c_4), .C(led_c_1), .Z(n18190)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_4_lut_then_3_lut.init = 16'h1010;
    LUT4 i1_4_lut_else_3_lut (.A(led_c_3), .B(led_c_0), .C(led_c_4), .D(led_c_1), 
         .Z(n18189)) /* synthesis lut_function=(!(A+(B (D)+!B (C+!(D))))) */ ;
    defparam i1_4_lut_else_3_lut.init = 16'h0144;
    LUT4 i2314_3_lut_4_lut (.A(n18138), .B(n18267), .C(led_c_3), .D(n187), 
         .Z(n12029)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2314_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_rep_164_3_lut_4_lut (.A(led_c_0), .B(n17963), .C(n26_adj_5659), 
         .D(led_c_4), .Z(n18134)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_2_lut_rep_164_3_lut_4_lut.init = 16'h0020;
    CCU2C _add_1_1436_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16700), .S0(cout_adj_5132));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1436_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1436_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_36 (.A0(d3_adj_5675[34]), .B0(d2_adj_5674[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[35]), .B1(d2_adj_5674[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16699), .COUT(n16700), .S0(d3_71__N_562_adj_5691[34]), 
          .S1(d3_71__N_562_adj_5691[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_34 (.A0(d3_adj_5675[32]), .B0(d2_adj_5674[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[33]), .B1(d2_adj_5674[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16698), .COUT(n16699), .S0(d3_71__N_562_adj_5691[32]), 
          .S1(d3_71__N_562_adj_5691[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_32 (.A0(d3_adj_5675[30]), .B0(d2_adj_5674[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[31]), .B1(d2_adj_5674[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16697), .COUT(n16698), .S0(d3_71__N_562_adj_5691[30]), 
          .S1(d3_71__N_562_adj_5691[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_30 (.A0(d3_adj_5675[28]), .B0(d2_adj_5674[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[29]), .B1(d2_adj_5674[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16696), .COUT(n16697), .S0(d3_71__N_562_adj_5691[28]), 
          .S1(d3_71__N_562_adj_5691[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_28 (.A0(d3_adj_5675[26]), .B0(d2_adj_5674[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[27]), .B1(d2_adj_5674[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16695), .COUT(n16696), .S0(d3_71__N_562_adj_5691[26]), 
          .S1(d3_71__N_562_adj_5691[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_26 (.A0(d3_adj_5675[24]), .B0(d2_adj_5674[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[25]), .B1(d2_adj_5674[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16694), .COUT(n16695), .S0(d3_71__N_562_adj_5691[24]), 
          .S1(d3_71__N_562_adj_5691[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_24 (.A0(d3_adj_5675[22]), .B0(d2_adj_5674[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[23]), .B1(d2_adj_5674[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16693), .COUT(n16694), .S0(d3_71__N_562_adj_5691[22]), 
          .S1(d3_71__N_562_adj_5691[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_22 (.A0(d3_adj_5675[20]), .B0(d2_adj_5674[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[21]), .B1(d2_adj_5674[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16692), .COUT(n16693), .S0(d3_71__N_562_adj_5691[20]), 
          .S1(d3_71__N_562_adj_5691[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_20 (.A0(d3_adj_5675[18]), .B0(d2_adj_5674[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[19]), .B1(d2_adj_5674[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16691), .COUT(n16692), .S0(d3_71__N_562_adj_5691[18]), 
          .S1(d3_71__N_562_adj_5691[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_18 (.A0(d3_adj_5675[16]), .B0(d2_adj_5674[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[17]), .B1(d2_adj_5674[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16690), .COUT(n16691), .S0(d3_71__N_562_adj_5691[16]), 
          .S1(d3_71__N_562_adj_5691[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_16 (.A0(d3_adj_5675[14]), .B0(d2_adj_5674[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[15]), .B1(d2_adj_5674[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16689), .COUT(n16690), .S0(d3_71__N_562_adj_5691[14]), 
          .S1(d3_71__N_562_adj_5691[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_14 (.A0(d3_adj_5675[12]), .B0(d2_adj_5674[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[13]), .B1(d2_adj_5674[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16688), .COUT(n16689), .S0(d3_71__N_562_adj_5691[12]), 
          .S1(d3_71__N_562_adj_5691[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_12 (.A0(d3_adj_5675[10]), .B0(d2_adj_5674[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[11]), .B1(d2_adj_5674[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16687), .COUT(n16688), .S0(d3_71__N_562_adj_5691[10]), 
          .S1(d3_71__N_562_adj_5691[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_10 (.A0(d3_adj_5675[8]), .B0(d2_adj_5674[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[9]), .B1(d2_adj_5674[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16686), .COUT(n16687), .S0(d3_71__N_562_adj_5691[8]), 
          .S1(d3_71__N_562_adj_5691[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_8 (.A0(d3_adj_5675[6]), .B0(d2_adj_5674[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[7]), .B1(d2_adj_5674[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16685), .COUT(n16686), .S0(d3_71__N_562_adj_5691[6]), 
          .S1(d3_71__N_562_adj_5691[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_6 (.A0(d3_adj_5675[4]), .B0(d2_adj_5674[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[5]), .B1(d2_adj_5674[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16684), .COUT(n16685), .S0(d3_71__N_562_adj_5691[4]), 
          .S1(d3_71__N_562_adj_5691[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_4 (.A0(d3_adj_5675[2]), .B0(d2_adj_5674[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[3]), .B1(d2_adj_5674[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16683), .COUT(n16684), .S0(d3_71__N_562_adj_5691[2]), 
          .S1(d3_71__N_562_adj_5691[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_2 (.A0(d3_adj_5675[0]), .B0(d2_adj_5674[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[1]), .B1(d2_adj_5674[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16683), .S1(d3_71__N_562_adj_5691[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1436_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_38 (.A0(d_d6_adj_5679[71]), .B0(d6_adj_5678[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16681), .S0(n78_adj_5354));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1628_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_36 (.A0(d_d6_adj_5679[69]), .B0(d6_adj_5678[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[70]), .B1(d6_adj_5678[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16680), .COUT(n16681), .S0(n84_adj_5356), 
          .S1(n81_adj_5355));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_34 (.A0(d_d6_adj_5679[67]), .B0(d6_adj_5678[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[68]), .B1(d6_adj_5678[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16679), .COUT(n16680), .S0(n90_adj_5358), 
          .S1(n87_adj_5357));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_32 (.A0(d_d6_adj_5679[65]), .B0(d6_adj_5678[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[66]), .B1(d6_adj_5678[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16678), .COUT(n16679), .S0(n96_adj_5360), 
          .S1(n93_adj_5359));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_30 (.A0(d_d6_adj_5679[63]), .B0(d6_adj_5678[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[64]), .B1(d6_adj_5678[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16677), .COUT(n16678), .S0(n102_adj_5362), 
          .S1(n99_adj_5361));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_30.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n317), .SP(clk_80mhz_enable_831), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n314), .SP(clk_80mhz_enable_831), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i4 (.D(n311), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n308), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i6 (.D(n305), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n302), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i8 (.D(n299), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i9 (.D(n296), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i10 (.D(n293), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n290), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i12 (.D(n287), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i13 (.D(n284), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i14 (.D(n281), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n278), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i16 (.D(n275), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i17 (.D(n272), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i18 (.D(n269), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n266), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i20 (.D(n263), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n260), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i22 (.D(n257), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i23 (.D(n254), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n251), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i25 (.D(n248), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n245), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i27 (.D(n242), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i28 (.D(n239), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i29 (.D(n236), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n233), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i31 (.D(n230), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n227), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i33 (.D(n224), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n221), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i35 (.D(n218), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i36 (.D(n215), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[36]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i37 (.D(n212), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i38 (.D(n209_adj_4996), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[38]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i39 (.D(n206), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i40 (.D(n203), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[40]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n200), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n197), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[42]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n194), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n191), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[44]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i45 (.D(n188), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i46 (.D(n185), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[46]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n182), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i48 (.D(n179), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[48]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i49 (.D(n176), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i50 (.D(n173), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[50]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i51 (.D(n170), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n167), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[52]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i53 (.D(n164), .SP(clk_80mhz_enable_881), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i54 (.D(n161), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[54]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i55 (.D(n158), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i56 (.D(n155), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[56]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n152), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i58 (.D(n149), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[58]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n146), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n143), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[60]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n140), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n137), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[62]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n134), .SP(clk_80mhz_enable_891), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    FD1P3AX CICGain__i2 (.D(led_c_1), .SP(clk_80mhz_enable_1470), .CK(clk_80mhz), 
            .Q(CICGain[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam CICGain__i2.GSR = "ENABLED";
    CCU2C _add_1_1628_add_4_28 (.A0(d_d6_adj_5679[61]), .B0(d6_adj_5678[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[62]), .B1(d6_adj_5678[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16676), .COUT(n16677), .S0(n108_adj_5364), 
          .S1(n105_adj_5363));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_6 (.A0(d_d9_adj_5685[39]), .B0(d9_adj_5684[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[40]), .B1(d9_adj_5684[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16496), .COUT(n16497));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_38 (.A0(d_d7[35]), .B0(d7[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16240), .S0(d8_71__N_1603[35]), .S1(cout_adj_5050));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1592_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_35 (.A0(d2_adj_5674[68]), .B0(cout_adj_5132), 
          .C0(n87_adj_5626), .D0(d3_adj_5675[68]), .A1(d2_adj_5674[69]), 
          .B1(cout_adj_5132), .C1(n84_adj_5625), .D1(d3_adj_5675[69]), 
          .CIN(n16052), .COUT(n16053), .S0(d3_71__N_562_adj_5691[68]), 
          .S1(d3_71__N_562_adj_5691[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_33 (.A0(d2_adj_5674[66]), .B0(cout_adj_5132), 
          .C0(n93_adj_5628), .D0(d3_adj_5675[66]), .A1(d2_adj_5674[67]), 
          .B1(cout_adj_5132), .C1(n90_adj_5627), .D1(d3_adj_5675[67]), 
          .CIN(n16051), .COUT(n16052), .S0(d3_71__N_562_adj_5691[66]), 
          .S1(d3_71__N_562_adj_5691[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_31 (.A0(d2_adj_5674[64]), .B0(cout_adj_5132), 
          .C0(n99_adj_5630), .D0(d3_adj_5675[64]), .A1(d2_adj_5674[65]), 
          .B1(cout_adj_5132), .C1(n96_adj_5629), .D1(d3_adj_5675[65]), 
          .CIN(n16050), .COUT(n16051), .S0(d3_71__N_562_adj_5691[64]), 
          .S1(d3_71__N_562_adj_5691[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_29 (.A0(d2_adj_5674[62]), .B0(cout_adj_5132), 
          .C0(n105_adj_5632), .D0(d3_adj_5675[62]), .A1(d2_adj_5674[63]), 
          .B1(cout_adj_5132), .C1(n102_adj_5631), .D1(d3_adj_5675[63]), 
          .CIN(n16049), .COUT(n16050), .S0(d3_71__N_562_adj_5691[62]), 
          .S1(d3_71__N_562_adj_5691[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_27 (.A0(d2_adj_5674[60]), .B0(cout_adj_5132), 
          .C0(n111_adj_5634), .D0(d3_adj_5675[60]), .A1(d2_adj_5674[61]), 
          .B1(cout_adj_5132), .C1(n108_adj_5633), .D1(d3_adj_5675[61]), 
          .CIN(n16048), .COUT(n16049), .S0(d3_71__N_562_adj_5691[60]), 
          .S1(d3_71__N_562_adj_5691[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_25 (.A0(d2_adj_5674[58]), .B0(cout_adj_5132), 
          .C0(n117_adj_5636), .D0(d3_adj_5675[58]), .A1(d2_adj_5674[59]), 
          .B1(cout_adj_5132), .C1(n114_adj_5635), .D1(d3_adj_5675[59]), 
          .CIN(n16047), .COUT(n16048), .S0(d3_71__N_562_adj_5691[58]), 
          .S1(d3_71__N_562_adj_5691[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_23 (.A0(d2_adj_5674[56]), .B0(cout_adj_5132), 
          .C0(n123_adj_5638), .D0(d3_adj_5675[56]), .A1(d2_adj_5674[57]), 
          .B1(cout_adj_5132), .C1(n120_adj_5637), .D1(d3_adj_5675[57]), 
          .CIN(n16046), .COUT(n16047), .S0(d3_71__N_562_adj_5691[56]), 
          .S1(d3_71__N_562_adj_5691[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_21 (.A0(d2_adj_5674[54]), .B0(cout_adj_5132), 
          .C0(n129_adj_5640), .D0(d3_adj_5675[54]), .A1(d2_adj_5674[55]), 
          .B1(cout_adj_5132), .C1(n126_adj_5639), .D1(d3_adj_5675[55]), 
          .CIN(n16045), .COUT(n16046), .S0(d3_71__N_562_adj_5691[54]), 
          .S1(d3_71__N_562_adj_5691[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_19 (.A0(d2_adj_5674[52]), .B0(cout_adj_5132), 
          .C0(n135_adj_5642), .D0(d3_adj_5675[52]), .A1(d2_adj_5674[53]), 
          .B1(cout_adj_5132), .C1(n132_adj_5641), .D1(d3_adj_5675[53]), 
          .CIN(n16044), .COUT(n16045), .S0(d3_71__N_562_adj_5691[52]), 
          .S1(d3_71__N_562_adj_5691[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_17 (.A0(d2_adj_5674[50]), .B0(cout_adj_5132), 
          .C0(n141_adj_5644), .D0(d3_adj_5675[50]), .A1(d2_adj_5674[51]), 
          .B1(cout_adj_5132), .C1(n138_adj_5643), .D1(d3_adj_5675[51]), 
          .CIN(n16043), .COUT(n16044), .S0(d3_71__N_562_adj_5691[50]), 
          .S1(d3_71__N_562_adj_5691[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_15 (.A0(d2_adj_5674[48]), .B0(cout_adj_5132), 
          .C0(n147_adj_5646), .D0(d3_adj_5675[48]), .A1(d2_adj_5674[49]), 
          .B1(cout_adj_5132), .C1(n144_adj_5645), .D1(d3_adj_5675[49]), 
          .CIN(n16042), .COUT(n16043), .S0(d3_71__N_562_adj_5691[48]), 
          .S1(d3_71__N_562_adj_5691[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_13 (.A0(d2_adj_5674[46]), .B0(cout_adj_5132), 
          .C0(n153_adj_5648), .D0(d3_adj_5675[46]), .A1(d2_adj_5674[47]), 
          .B1(cout_adj_5132), .C1(n150_adj_5647), .D1(d3_adj_5675[47]), 
          .CIN(n16041), .COUT(n16042), .S0(d3_71__N_562_adj_5691[46]), 
          .S1(d3_71__N_562_adj_5691[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_11 (.A0(d2_adj_5674[44]), .B0(cout_adj_5132), 
          .C0(n159_adj_5650), .D0(d3_adj_5675[44]), .A1(d2_adj_5674[45]), 
          .B1(cout_adj_5132), .C1(n156_adj_5649), .D1(d3_adj_5675[45]), 
          .CIN(n16040), .COUT(n16041), .S0(d3_71__N_562_adj_5691[44]), 
          .S1(d3_71__N_562_adj_5691[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_9 (.A0(d2_adj_5674[42]), .B0(cout_adj_5132), 
          .C0(n165_adj_5652), .D0(d3_adj_5675[42]), .A1(d2_adj_5674[43]), 
          .B1(cout_adj_5132), .C1(n162_adj_5651), .D1(d3_adj_5675[43]), 
          .CIN(n16039), .COUT(n16040), .S0(d3_71__N_562_adj_5691[42]), 
          .S1(d3_71__N_562_adj_5691[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_7 (.A0(d2_adj_5674[40]), .B0(cout_adj_5132), 
          .C0(n171_adj_5654), .D0(d3_adj_5675[40]), .A1(d2_adj_5674[41]), 
          .B1(cout_adj_5132), .C1(n168_adj_5653), .D1(d3_adj_5675[41]), 
          .CIN(n16038), .COUT(n16039), .S0(d3_71__N_562_adj_5691[40]), 
          .S1(d3_71__N_562_adj_5691[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_5 (.A0(d2_adj_5674[38]), .B0(cout_adj_5132), 
          .C0(n177_adj_5656), .D0(d3_adj_5675[38]), .A1(d2_adj_5674[39]), 
          .B1(cout_adj_5132), .C1(n174_adj_5655), .D1(d3_adj_5675[39]), 
          .CIN(n16037), .COUT(n16038), .S0(d3_71__N_562_adj_5691[38]), 
          .S1(d3_71__N_562_adj_5691[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_3 (.A0(d2_adj_5674[36]), .B0(cout_adj_5132), 
          .C0(n183_adj_5658), .D0(d3_adj_5675[36]), .A1(d2_adj_5674[37]), 
          .B1(cout_adj_5132), .C1(n180_adj_5657), .D1(d3_adj_5675[37]), 
          .CIN(n16036), .COUT(n16037), .S0(d3_71__N_562_adj_5691[36]), 
          .S1(d3_71__N_562_adj_5691[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5132), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16036));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1496_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1496_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_37 (.A0(d1_adj_5673[70]), .B0(cout_adj_5131), 
          .C0(n81_adj_2805), .D0(d2_adj_5674[70]), .A1(d1_adj_5673[71]), 
          .B1(cout_adj_5131), .C1(n78_adj_2806), .D1(d2_adj_5674[71]), 
          .CIN(n16031), .S0(d2_71__N_490_adj_5690[70]), .S1(d2_71__N_490_adj_5690[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_35 (.A0(d1_adj_5673[68]), .B0(cout_adj_5131), 
          .C0(n87_adj_2803), .D0(d2_adj_5674[68]), .A1(d1_adj_5673[69]), 
          .B1(cout_adj_5131), .C1(n84_adj_2804), .D1(d2_adj_5674[69]), 
          .CIN(n16030), .COUT(n16031), .S0(d2_71__N_490_adj_5690[68]), 
          .S1(d2_71__N_490_adj_5690[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_33 (.A0(d1_adj_5673[66]), .B0(cout_adj_5131), 
          .C0(n93_adj_2801), .D0(d2_adj_5674[66]), .A1(d1_adj_5673[67]), 
          .B1(cout_adj_5131), .C1(n90_adj_2802), .D1(d2_adj_5674[67]), 
          .CIN(n16029), .COUT(n16030), .S0(d2_71__N_490_adj_5690[66]), 
          .S1(d2_71__N_490_adj_5690[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_31 (.A0(d1_adj_5673[64]), .B0(cout_adj_5131), 
          .C0(n99_adj_2799), .D0(d2_adj_5674[64]), .A1(d1_adj_5673[65]), 
          .B1(cout_adj_5131), .C1(n96_adj_2800), .D1(d2_adj_5674[65]), 
          .CIN(n16028), .COUT(n16029), .S0(d2_71__N_490_adj_5690[64]), 
          .S1(d2_71__N_490_adj_5690[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_29 (.A0(d1_adj_5673[62]), .B0(cout_adj_5131), 
          .C0(n105_adj_2797), .D0(d2_adj_5674[62]), .A1(d1_adj_5673[63]), 
          .B1(cout_adj_5131), .C1(n102_adj_2798), .D1(d2_adj_5674[63]), 
          .CIN(n16027), .COUT(n16028), .S0(d2_71__N_490_adj_5690[62]), 
          .S1(d2_71__N_490_adj_5690[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_27 (.A0(d1_adj_5673[60]), .B0(cout_adj_5131), 
          .C0(n111_adj_2795), .D0(d2_adj_5674[60]), .A1(d1_adj_5673[61]), 
          .B1(cout_adj_5131), .C1(n108_adj_2796), .D1(d2_adj_5674[61]), 
          .CIN(n16026), .COUT(n16027), .S0(d2_71__N_490_adj_5690[60]), 
          .S1(d2_71__N_490_adj_5690[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_25 (.A0(d1_adj_5673[58]), .B0(cout_adj_5131), 
          .C0(n117_adj_2793), .D0(d2_adj_5674[58]), .A1(d1_adj_5673[59]), 
          .B1(cout_adj_5131), .C1(n114_adj_2794), .D1(d2_adj_5674[59]), 
          .CIN(n16025), .COUT(n16026), .S0(d2_71__N_490_adj_5690[58]), 
          .S1(d2_71__N_490_adj_5690[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_23 (.A0(d1_adj_5673[56]), .B0(cout_adj_5131), 
          .C0(n123_adj_2791), .D0(d2_adj_5674[56]), .A1(d1_adj_5673[57]), 
          .B1(cout_adj_5131), .C1(n120_adj_2792), .D1(d2_adj_5674[57]), 
          .CIN(n16024), .COUT(n16025), .S0(d2_71__N_490_adj_5690[56]), 
          .S1(d2_71__N_490_adj_5690[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_21 (.A0(d1_adj_5673[54]), .B0(cout_adj_5131), 
          .C0(n129_adj_2789), .D0(d2_adj_5674[54]), .A1(d1_adj_5673[55]), 
          .B1(cout_adj_5131), .C1(n126_adj_2790), .D1(d2_adj_5674[55]), 
          .CIN(n16023), .COUT(n16024), .S0(d2_71__N_490_adj_5690[54]), 
          .S1(d2_71__N_490_adj_5690[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_19 (.A0(d1_adj_5673[52]), .B0(cout_adj_5131), 
          .C0(n135_adj_2787), .D0(d2_adj_5674[52]), .A1(d1_adj_5673[53]), 
          .B1(cout_adj_5131), .C1(n132_adj_2788), .D1(d2_adj_5674[53]), 
          .CIN(n16022), .COUT(n16023), .S0(d2_71__N_490_adj_5690[52]), 
          .S1(d2_71__N_490_adj_5690[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_17 (.A0(d1_adj_5673[50]), .B0(cout_adj_5131), 
          .C0(n141_adj_2785), .D0(d2_adj_5674[50]), .A1(d1_adj_5673[51]), 
          .B1(cout_adj_5131), .C1(n138_adj_2786), .D1(d2_adj_5674[51]), 
          .CIN(n16021), .COUT(n16022), .S0(d2_71__N_490_adj_5690[50]), 
          .S1(d2_71__N_490_adj_5690[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_15 (.A0(d1_adj_5673[48]), .B0(cout_adj_5131), 
          .C0(n147_adj_2783), .D0(d2_adj_5674[48]), .A1(d1_adj_5673[49]), 
          .B1(cout_adj_5131), .C1(n144_adj_2784), .D1(d2_adj_5674[49]), 
          .CIN(n16020), .COUT(n16021), .S0(d2_71__N_490_adj_5690[48]), 
          .S1(d2_71__N_490_adj_5690[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_13 (.A0(d1_adj_5673[46]), .B0(cout_adj_5131), 
          .C0(n153_adj_2781), .D0(d2_adj_5674[46]), .A1(d1_adj_5673[47]), 
          .B1(cout_adj_5131), .C1(n150_adj_2782), .D1(d2_adj_5674[47]), 
          .CIN(n16019), .COUT(n16020), .S0(d2_71__N_490_adj_5690[46]), 
          .S1(d2_71__N_490_adj_5690[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_11 (.A0(d1_adj_5673[44]), .B0(cout_adj_5131), 
          .C0(n159_adj_2779), .D0(d2_adj_5674[44]), .A1(d1_adj_5673[45]), 
          .B1(cout_adj_5131), .C1(n156_adj_2780), .D1(d2_adj_5674[45]), 
          .CIN(n16018), .COUT(n16019), .S0(d2_71__N_490_adj_5690[44]), 
          .S1(d2_71__N_490_adj_5690[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_9 (.A0(d1_adj_5673[42]), .B0(cout_adj_5131), 
          .C0(n165_adj_2777), .D0(d2_adj_5674[42]), .A1(d1_adj_5673[43]), 
          .B1(cout_adj_5131), .C1(n162_adj_2778), .D1(d2_adj_5674[43]), 
          .CIN(n16017), .COUT(n16018), .S0(d2_71__N_490_adj_5690[42]), 
          .S1(d2_71__N_490_adj_5690[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_7 (.A0(d1_adj_5673[40]), .B0(cout_adj_5131), 
          .C0(n171_adj_2775), .D0(d2_adj_5674[40]), .A1(d1_adj_5673[41]), 
          .B1(cout_adj_5131), .C1(n168_adj_2776), .D1(d2_adj_5674[41]), 
          .CIN(n16016), .COUT(n16017), .S0(d2_71__N_490_adj_5690[40]), 
          .S1(d2_71__N_490_adj_5690[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_5 (.A0(d1_adj_5673[38]), .B0(cout_adj_5131), 
          .C0(n177_adj_2773), .D0(d2_adj_5674[38]), .A1(d1_adj_5673[39]), 
          .B1(cout_adj_5131), .C1(n174_adj_2774), .D1(d2_adj_5674[39]), 
          .CIN(n16015), .COUT(n16016), .S0(d2_71__N_490_adj_5690[38]), 
          .S1(d2_71__N_490_adj_5690[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_3 (.A0(d1_adj_5673[36]), .B0(cout_adj_5131), 
          .C0(n183_adj_2771), .D0(d2_adj_5674[36]), .A1(d1_adj_5673[37]), 
          .B1(cout_adj_5131), .C1(n180_adj_2772), .D1(d2_adj_5674[37]), 
          .CIN(n16014), .COUT(n16015), .S0(d2_71__N_490_adj_5690[36]), 
          .S1(d2_71__N_490_adj_5690[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5131), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16014));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1499_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1499_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_38 (.A0(d2_adj_5674[71]), .B0(d1_adj_5673[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16010), .S0(n78_adj_2806));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1571_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_36 (.A0(d2_adj_5674[69]), .B0(d1_adj_5673[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[70]), .B1(d1_adj_5673[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16009), .COUT(n16010), .S0(n84_adj_2804), 
          .S1(n81_adj_2805));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_34 (.A0(d2_adj_5674[67]), .B0(d1_adj_5673[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[68]), .B1(d1_adj_5673[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16008), .COUT(n16009), .S0(n90_adj_2802), 
          .S1(n87_adj_2803));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_32 (.A0(d2_adj_5674[65]), .B0(d1_adj_5673[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[66]), .B1(d1_adj_5673[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16007), .COUT(n16008), .S0(n96_adj_2800), 
          .S1(n93_adj_2801));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_30 (.A0(d2_adj_5674[63]), .B0(d1_adj_5673[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[64]), .B1(d1_adj_5673[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16006), .COUT(n16007), .S0(n102_adj_2798), 
          .S1(n99_adj_2799));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_28 (.A0(d2_adj_5674[61]), .B0(d1_adj_5673[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[62]), .B1(d1_adj_5673[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16005), .COUT(n16006), .S0(n108_adj_2796), 
          .S1(n105_adj_2797));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_26 (.A0(d2_adj_5674[59]), .B0(d1_adj_5673[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[60]), .B1(d1_adj_5673[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16004), .COUT(n16005), .S0(n114_adj_2794), 
          .S1(n111_adj_2795));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_24 (.A0(d2_adj_5674[57]), .B0(d1_adj_5673[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[58]), .B1(d1_adj_5673[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16003), .COUT(n16004), .S0(n120_adj_2792), 
          .S1(n117_adj_2793));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_22 (.A0(d2_adj_5674[55]), .B0(d1_adj_5673[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[56]), .B1(d1_adj_5673[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16002), .COUT(n16003), .S0(n126_adj_2790), 
          .S1(n123_adj_2791));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_20 (.A0(d2_adj_5674[53]), .B0(d1_adj_5673[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[54]), .B1(d1_adj_5673[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16001), .COUT(n16002), .S0(n132_adj_2788), 
          .S1(n129_adj_2789));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_18 (.A0(d2_adj_5674[51]), .B0(d1_adj_5673[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[52]), .B1(d1_adj_5673[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16000), .COUT(n16001), .S0(n138_adj_2786), 
          .S1(n135_adj_2787));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_16 (.A0(d2_adj_5674[49]), .B0(d1_adj_5673[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[50]), .B1(d1_adj_5673[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15999), .COUT(n16000), .S0(n144_adj_2784), 
          .S1(n141_adj_2785));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_14 (.A0(d2_adj_5674[47]), .B0(d1_adj_5673[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[48]), .B1(d1_adj_5673[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15998), .COUT(n15999), .S0(n150_adj_2782), 
          .S1(n147_adj_2783));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_12 (.A0(d2_adj_5674[45]), .B0(d1_adj_5673[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[46]), .B1(d1_adj_5673[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15997), .COUT(n15998), .S0(n156_adj_2780), 
          .S1(n153_adj_2781));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_10 (.A0(d2_adj_5674[43]), .B0(d1_adj_5673[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[44]), .B1(d1_adj_5673[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15996), .COUT(n15997), .S0(n162_adj_2778), 
          .S1(n159_adj_2779));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_8 (.A0(d2_adj_5674[41]), .B0(d1_adj_5673[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[42]), .B1(d1_adj_5673[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15995), .COUT(n15996), .S0(n168_adj_2776), 
          .S1(n165_adj_2777));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_6 (.A0(d2_adj_5674[39]), .B0(d1_adj_5673[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[40]), .B1(d1_adj_5673[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15994), .COUT(n15995), .S0(n174_adj_2774), 
          .S1(n171_adj_2775));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_4 (.A0(d2_adj_5674[37]), .B0(d1_adj_5673[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[38]), .B1(d1_adj_5673[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15993), .COUT(n15994), .S0(n180_adj_2772), 
          .S1(n177_adj_2773));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2_adj_5674[36]), .B1(d1_adj_5673[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15993), .S1(n183_adj_2771));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1571_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1571_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_38 (.A0(d_d6[35]), .B0(d6[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15992), .S0(d7_71__N_1531[35]), .S1(cout_adj_5490));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1523_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_36 (.A0(d_d6[33]), .B0(d6[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[34]), .B1(d6[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15991), .COUT(n15992), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_34 (.A0(d_d6[31]), .B0(d6[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[32]), .B1(d6[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15990), .COUT(n15991), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_32 (.A0(d_d6[29]), .B0(d6[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[30]), .B1(d6[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15989), .COUT(n15990), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_26 (.A0(d_d6_adj_5679[59]), .B0(d6_adj_5678[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[60]), .B1(d6_adj_5678[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16675), .COUT(n16676), .S0(n114_adj_5366), 
          .S1(n111_adj_5365));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_24 (.A0(d_d6_adj_5679[57]), .B0(d6_adj_5678[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[58]), .B1(d6_adj_5678[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16674), .COUT(n16675), .S0(n120_adj_5368), 
          .S1(n117_adj_5367));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_22 (.A0(d_d6_adj_5679[55]), .B0(d6_adj_5678[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[56]), .B1(d6_adj_5678[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16673), .COUT(n16674), .S0(n126_adj_5370), 
          .S1(n123_adj_5369));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_20 (.A0(d_d6_adj_5679[53]), .B0(d6_adj_5678[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[54]), .B1(d6_adj_5678[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16672), .COUT(n16673), .S0(n132_adj_5372), 
          .S1(n129_adj_5371));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_18 (.A0(d_d6_adj_5679[51]), .B0(d6_adj_5678[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[52]), .B1(d6_adj_5678[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16671), .COUT(n16672), .S0(n138_adj_5374), 
          .S1(n135_adj_5373));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_16 (.A0(d_d6_adj_5679[49]), .B0(d6_adj_5678[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[50]), .B1(d6_adj_5678[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16670), .COUT(n16671), .S0(n144_adj_5376), 
          .S1(n141_adj_5375));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_14 (.A0(d_d6_adj_5679[47]), .B0(d6_adj_5678[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[48]), .B1(d6_adj_5678[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16669), .COUT(n16670), .S0(n150_adj_5378), 
          .S1(n147_adj_5377));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_12 (.A0(d_d6_adj_5679[45]), .B0(d6_adj_5678[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[46]), .B1(d6_adj_5678[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16668), .COUT(n16669), .S0(n156_adj_5380), 
          .S1(n153_adj_5379));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_10 (.A0(d_d6_adj_5679[43]), .B0(d6_adj_5678[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[44]), .B1(d6_adj_5678[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16667), .COUT(n16668), .S0(n162_adj_5382), 
          .S1(n159_adj_5381));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_31 (.A0(d_tmp[64]), .B0(cout_adj_5496), .C0(n99_adj_5058), 
          .D0(n9_adj_4761), .A1(d_tmp[65]), .B1(cout_adj_5496), .C1(n96_adj_5057), 
          .D1(n8_adj_4762), .CIN(n16338), .COUT(n16339), .S0(d6_71__N_1459[64]), 
          .S1(d6_71__N_1459[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_8 (.A0(d_d6_adj_5679[41]), .B0(d6_adj_5678[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[42]), .B1(d6_adj_5678[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16666), .COUT(n16667), .S0(n168_adj_5384), 
          .S1(n165_adj_5383));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4998), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16368));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1487_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1487_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_24 (.A0(d4_adj_5676[57]), .B0(d3_adj_5675[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[58]), .B1(d3_adj_5675[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16278), .COUT(n16279), .S0(n120_adj_4746), 
          .S1(n117_adj_4745));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_6 (.A0(d_d6_adj_5679[39]), .B0(d6_adj_5678[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[40]), .B1(d6_adj_5678[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16665), .COUT(n16666), .S0(n174_adj_5386), 
          .S1(n171_adj_5385));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_22 (.A0(d4_adj_5676[55]), .B0(d3_adj_5675[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[56]), .B1(d3_adj_5675[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16277), .COUT(n16278), .S0(n126_adj_4788), 
          .S1(n123_adj_4747));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_4 (.A0(d_d9_adj_5685[37]), .B0(d9_adj_5684[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[38]), .B1(d9_adj_5684[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16495), .COUT(n16496));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_4.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_171_4_lut (.A(led_c_0), .B(n17963), .C(led_c_4), 
         .D(n26_adj_5659), .Z(n18141)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_3_lut_rep_171_4_lut.init = 16'h2000;
    CCU2C _add_1_1577_add_4_20 (.A0(d4_adj_5676[53]), .B0(d3_adj_5675[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[54]), .B1(d3_adj_5675[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16276), .COUT(n16277), .S0(n132_adj_4790), 
          .S1(n129_adj_4789));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_36 (.A0(d_d7[33]), .B0(d7[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[34]), .B1(d7[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16239), .COUT(n16240), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_34 (.A0(d_d7[31]), .B0(d7[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[32]), .B1(d7[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16238), .COUT(n16239), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_32 (.A0(d_d7[29]), .B0(d7[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[30]), .B1(d7[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16237), .COUT(n16238), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_30 (.A0(d_d6[27]), .B0(d6[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[28]), .B1(d6[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15988), .COUT(n15989), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_28 (.A0(d_d6[25]), .B0(d6[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[26]), .B1(d6[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15987), .COUT(n15988), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_26 (.A0(d_d6[23]), .B0(d6[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[24]), .B1(d6[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15986), .COUT(n15987), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_24 (.A0(d_d6[21]), .B0(d6[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[22]), .B1(d6[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15985), .COUT(n15986), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_22 (.A0(d_d6[19]), .B0(d6[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[20]), .B1(d6[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15984), .COUT(n15985), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_20 (.A0(d_d6[17]), .B0(d6[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[18]), .B1(d6[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15983), .COUT(n15984), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_18 (.A0(d_d6[15]), .B0(d6[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[16]), .B1(d6[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15982), .COUT(n15983), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_16 (.A0(d_d6[13]), .B0(d6[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[14]), .B1(d6[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15981), .COUT(n15982), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_14 (.A0(d_d6[11]), .B0(d6[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[12]), .B1(d6[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15980), .COUT(n15981), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_12 (.A0(d_d6[9]), .B0(d6[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[10]), .B1(d6[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15979), .COUT(n15980), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_10 (.A0(d_d6[7]), .B0(d6[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[8]), .B1(d6[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15978), .COUT(n15979), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_8 (.A0(d_d6[5]), .B0(d6[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[6]), .B1(d6[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15977), .COUT(n15978), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_6 (.A0(d_d6[3]), .B0(d6[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[4]), .B1(d6[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15976), .COUT(n15977), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_4 (.A0(d_d6[1]), .B0(d6[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[2]), .B1(d6[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15975), .COUT(n15976), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[0]), .B1(d6[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15975), .S1(d7_71__N_1531[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1523_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_38 (.A0(d_d6_adj_5679[35]), .B0(d6_adj_5678[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15974), .S0(d7_71__N_1531_adj_5706[35]), 
          .S1(cout_adj_5192));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1607_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_36 (.A0(d_d6_adj_5679[33]), .B0(d6_adj_5678[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[34]), .B1(d6_adj_5678[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15973), .COUT(n15974), .S0(d7_71__N_1531_adj_5706[33]), 
          .S1(d7_71__N_1531_adj_5706[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_34 (.A0(d_d6_adj_5679[31]), .B0(d6_adj_5678[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[32]), .B1(d6_adj_5678[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15972), .COUT(n15973), .S0(d7_71__N_1531_adj_5706[31]), 
          .S1(d7_71__N_1531_adj_5706[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_32 (.A0(d_d6_adj_5679[29]), .B0(d6_adj_5678[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[30]), .B1(d6_adj_5678[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15971), .COUT(n15972), .S0(d7_71__N_1531_adj_5706[29]), 
          .S1(d7_71__N_1531_adj_5706[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_30 (.A0(d_d6_adj_5679[27]), .B0(d6_adj_5678[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[28]), .B1(d6_adj_5678[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15970), .COUT(n15971), .S0(d7_71__N_1531_adj_5706[27]), 
          .S1(d7_71__N_1531_adj_5706[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_28 (.A0(d_d6_adj_5679[25]), .B0(d6_adj_5678[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[26]), .B1(d6_adj_5678[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15969), .COUT(n15970), .S0(d7_71__N_1531_adj_5706[25]), 
          .S1(d7_71__N_1531_adj_5706[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_26 (.A0(d_d6_adj_5679[23]), .B0(d6_adj_5678[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[24]), .B1(d6_adj_5678[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15968), .COUT(n15969), .S0(d7_71__N_1531_adj_5706[23]), 
          .S1(d7_71__N_1531_adj_5706[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_24 (.A0(d_d6_adj_5679[21]), .B0(d6_adj_5678[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[22]), .B1(d6_adj_5678[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15967), .COUT(n15968), .S0(d7_71__N_1531_adj_5706[21]), 
          .S1(d7_71__N_1531_adj_5706[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_22 (.A0(d_d6_adj_5679[19]), .B0(d6_adj_5678[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[20]), .B1(d6_adj_5678[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15966), .COUT(n15967), .S0(d7_71__N_1531_adj_5706[19]), 
          .S1(d7_71__N_1531_adj_5706[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_20 (.A0(d_d6_adj_5679[17]), .B0(d6_adj_5678[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[18]), .B1(d6_adj_5678[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15965), .COUT(n15966), .S0(d7_71__N_1531_adj_5706[17]), 
          .S1(d7_71__N_1531_adj_5706[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_18 (.A0(d_d6_adj_5679[15]), .B0(d6_adj_5678[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[16]), .B1(d6_adj_5678[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15964), .COUT(n15965), .S0(d7_71__N_1531_adj_5706[15]), 
          .S1(d7_71__N_1531_adj_5706[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_16 (.A0(d_d6_adj_5679[13]), .B0(d6_adj_5678[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[14]), .B1(d6_adj_5678[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15963), .COUT(n15964), .S0(d7_71__N_1531_adj_5706[13]), 
          .S1(d7_71__N_1531_adj_5706[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_14 (.A0(d_d6_adj_5679[11]), .B0(d6_adj_5678[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[12]), .B1(d6_adj_5678[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15962), .COUT(n15963), .S0(d7_71__N_1531_adj_5706[11]), 
          .S1(d7_71__N_1531_adj_5706[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_12 (.A0(d_d6_adj_5679[9]), .B0(d6_adj_5678[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[10]), .B1(d6_adj_5678[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15961), .COUT(n15962), .S0(d7_71__N_1531_adj_5706[9]), 
          .S1(d7_71__N_1531_adj_5706[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_10 (.A0(d_d6_adj_5679[7]), .B0(d6_adj_5678[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[8]), .B1(d6_adj_5678[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15960), .COUT(n15961), .S0(d7_71__N_1531_adj_5706[7]), 
          .S1(d7_71__N_1531_adj_5706[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_8 (.A0(d_d6_adj_5679[5]), .B0(d6_adj_5678[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[6]), .B1(d6_adj_5678[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15959), .COUT(n15960), .S0(d7_71__N_1531_adj_5706[5]), 
          .S1(d7_71__N_1531_adj_5706[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_6 (.A0(d_d6_adj_5679[3]), .B0(d6_adj_5678[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[4]), .B1(d6_adj_5678[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15958), .COUT(n15959), .S0(d7_71__N_1531_adj_5706[3]), 
          .S1(d7_71__N_1531_adj_5706[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_4 (.A0(d_d6_adj_5679[1]), .B0(d6_adj_5678[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[2]), .B1(d6_adj_5678[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15957), .COUT(n15958), .S0(d7_71__N_1531_adj_5706[1]), 
          .S1(d7_71__N_1531_adj_5706[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1607_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5679[0]), .B1(d6_adj_5678[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15957), .S1(d7_71__N_1531_adj_5706[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1607_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1607_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1607_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_37 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n81_adj_5577), .D0(d1_adj_5673[70]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n78_adj_5576), .D1(d1_adj_5673[71]), 
          .CIN(n15955), .S0(d1_71__N_418_adj_5689[70]), .S1(d1_71__N_418_adj_5689[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_35 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n87_adj_5579), .D0(d1_adj_5673[68]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n84_adj_5578), .D1(d1_adj_5673[69]), 
          .CIN(n15954), .COUT(n15955), .S0(d1_71__N_418_adj_5689[68]), 
          .S1(d1_71__N_418_adj_5689[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_33 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n93_adj_5581), .D0(d1_adj_5673[66]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n90_adj_5580), .D1(d1_adj_5673[67]), 
          .CIN(n15953), .COUT(n15954), .S0(d1_71__N_418_adj_5689[66]), 
          .S1(d1_71__N_418_adj_5689[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_31 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n99_adj_5583), .D0(d1_adj_5673[64]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n96_adj_5582), .D1(d1_adj_5673[65]), 
          .CIN(n15952), .COUT(n15953), .S0(d1_71__N_418_adj_5689[64]), 
          .S1(d1_71__N_418_adj_5689[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_29 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n105_adj_5585), .D0(d1_adj_5673[62]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n102_adj_5584), .D1(d1_adj_5673[63]), 
          .CIN(n15951), .COUT(n15952), .S0(d1_71__N_418_adj_5689[62]), 
          .S1(d1_71__N_418_adj_5689[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_27 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n111_adj_5587), .D0(d1_adj_5673[60]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n108_adj_5586), .D1(d1_adj_5673[61]), 
          .CIN(n15950), .COUT(n15951), .S0(d1_71__N_418_adj_5689[60]), 
          .S1(d1_71__N_418_adj_5689[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_25 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n117_adj_5589), .D0(d1_adj_5673[58]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n114_adj_5588), .D1(d1_adj_5673[59]), 
          .CIN(n15949), .COUT(n15950), .S0(d1_71__N_418_adj_5689[58]), 
          .S1(d1_71__N_418_adj_5689[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_23 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n123_adj_5591), .D0(d1_adj_5673[56]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n120_adj_5590), .D1(d1_adj_5673[57]), 
          .CIN(n15948), .COUT(n15949), .S0(d1_71__N_418_adj_5689[56]), 
          .S1(d1_71__N_418_adj_5689[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_21 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n129_adj_5593), .D0(d1_adj_5673[54]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n126_adj_5592), .D1(d1_adj_5673[55]), 
          .CIN(n15947), .COUT(n15948), .S0(d1_71__N_418_adj_5689[54]), 
          .S1(d1_71__N_418_adj_5689[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_19 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n135_adj_5595), .D0(d1_adj_5673[52]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n132_adj_5594), .D1(d1_adj_5673[53]), 
          .CIN(n15946), .COUT(n15947), .S0(d1_71__N_418_adj_5689[52]), 
          .S1(d1_71__N_418_adj_5689[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_17 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n141_adj_5597), .D0(d1_adj_5673[50]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n138_adj_5596), .D1(d1_adj_5673[51]), 
          .CIN(n15945), .COUT(n15946), .S0(d1_71__N_418_adj_5689[50]), 
          .S1(d1_71__N_418_adj_5689[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_15 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n147_adj_5599), .D0(d1_adj_5673[48]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n144_adj_5598), .D1(d1_adj_5673[49]), 
          .CIN(n15944), .COUT(n15945), .S0(d1_71__N_418_adj_5689[48]), 
          .S1(d1_71__N_418_adj_5689[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_13 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n153_adj_5601), .D0(d1_adj_5673[46]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n150_adj_5600), .D1(d1_adj_5673[47]), 
          .CIN(n15943), .COUT(n15944), .S0(d1_71__N_418_adj_5689[46]), 
          .S1(d1_71__N_418_adj_5689[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_11 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n159_adj_5603), .D0(d1_adj_5673[44]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n156_adj_5602), .D1(d1_adj_5673[45]), 
          .CIN(n15942), .COUT(n15943), .S0(d1_71__N_418_adj_5689[44]), 
          .S1(d1_71__N_418_adj_5689[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_9 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n165_adj_5605), .D0(d1_adj_5673[42]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n162_adj_5604), .D1(d1_adj_5673[43]), 
          .CIN(n15941), .COUT(n15942), .S0(d1_71__N_418_adj_5689[42]), 
          .S1(d1_71__N_418_adj_5689[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_7 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n171_adj_5607), .D0(d1_adj_5673[40]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n168_adj_5606), .D1(d1_adj_5673[41]), 
          .CIN(n15940), .COUT(n15941), .S0(d1_71__N_418_adj_5689[40]), 
          .S1(d1_71__N_418_adj_5689[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_5 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n177_adj_5609), .D0(d1_adj_5673[38]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n174_adj_5608), .D1(d1_adj_5673[39]), 
          .CIN(n15939), .COUT(n15940), .S0(d1_71__N_418_adj_5689[38]), 
          .S1(d1_71__N_418_adj_5689[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_3 (.A0(MixerOutCos[11]), .B0(cout_adj_5089), 
          .C0(n183_adj_5611), .D0(d1_adj_5673[36]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5089), .C1(n180_adj_5610), .D1(d1_adj_5673[37]), 
          .CIN(n15938), .COUT(n15939), .S0(d1_71__N_418_adj_5689[36]), 
          .S1(d1_71__N_418_adj_5689[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5089), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15938));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1502_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1502_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_38 (.A0(d_d_tmp_adj_5672[71]), .B0(d_tmp_adj_5671[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15934), .S0(n78_adj_5318));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1625_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_36 (.A0(d_d_tmp_adj_5672[69]), .B0(d_tmp_adj_5671[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[70]), .B1(d_tmp_adj_5671[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15933), .COUT(n15934), .S0(n84_adj_5320), 
          .S1(n81_adj_5319));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_34 (.A0(d_d_tmp_adj_5672[67]), .B0(d_tmp_adj_5671[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[68]), .B1(d_tmp_adj_5671[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15932), .COUT(n15933), .S0(n90_adj_5322), 
          .S1(n87_adj_5321));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_32 (.A0(d_d_tmp_adj_5672[65]), .B0(d_tmp_adj_5671[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[66]), .B1(d_tmp_adj_5671[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15931), .COUT(n15932), .S0(n96_adj_5324), 
          .S1(n93_adj_5323));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_30 (.A0(d_d_tmp_adj_5672[63]), .B0(d_tmp_adj_5671[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[64]), .B1(d_tmp_adj_5671[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15930), .COUT(n15931), .S0(n102_adj_5326), 
          .S1(n99_adj_5325));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_28 (.A0(d_d_tmp_adj_5672[61]), .B0(d_tmp_adj_5671[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[62]), .B1(d_tmp_adj_5671[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15929), .COUT(n15930), .S0(n108_adj_5328), 
          .S1(n105_adj_5327));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_26 (.A0(d_d_tmp_adj_5672[59]), .B0(d_tmp_adj_5671[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[60]), .B1(d_tmp_adj_5671[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15928), .COUT(n15929), .S0(n114_adj_5330), 
          .S1(n111_adj_5329));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_24 (.A0(d_d_tmp_adj_5672[57]), .B0(d_tmp_adj_5671[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[58]), .B1(d_tmp_adj_5671[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15927), .COUT(n15928), .S0(n120_adj_5332), 
          .S1(n117_adj_5331));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_22 (.A0(d_d_tmp_adj_5672[55]), .B0(d_tmp_adj_5671[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[56]), .B1(d_tmp_adj_5671[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15926), .COUT(n15927), .S0(n126_adj_5334), 
          .S1(n123_adj_5333));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_20 (.A0(d_d_tmp_adj_5672[53]), .B0(d_tmp_adj_5671[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[54]), .B1(d_tmp_adj_5671[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15925), .COUT(n15926), .S0(n132_adj_5336), 
          .S1(n129_adj_5335));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_18 (.A0(d_d_tmp_adj_5672[51]), .B0(d_tmp_adj_5671[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[52]), .B1(d_tmp_adj_5671[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15924), .COUT(n15925), .S0(n138_adj_5338), 
          .S1(n135_adj_5337));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_16 (.A0(d_d_tmp_adj_5672[49]), .B0(d_tmp_adj_5671[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[50]), .B1(d_tmp_adj_5671[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15923), .COUT(n15924), .S0(n144_adj_5340), 
          .S1(n141_adj_5339));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_14 (.A0(d_d_tmp_adj_5672[47]), .B0(d_tmp_adj_5671[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[48]), .B1(d_tmp_adj_5671[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15922), .COUT(n15923), .S0(n150_adj_5342), 
          .S1(n147_adj_5341));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_12 (.A0(d_d_tmp_adj_5672[45]), .B0(d_tmp_adj_5671[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[46]), .B1(d_tmp_adj_5671[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15921), .COUT(n15922), .S0(n156_adj_5344), 
          .S1(n153_adj_5343));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_10 (.A0(d_d_tmp_adj_5672[43]), .B0(d_tmp_adj_5671[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[44]), .B1(d_tmp_adj_5671[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15920), .COUT(n15921), .S0(n162_adj_5346), 
          .S1(n159_adj_5345));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_10.INJECT1_1 = "NO";
    LUT4 i5643_2_lut (.A(MultResult2[0]), .B(MultResult1[0]), .Z(n126_adj_5191)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5643_2_lut.init = 16'h6666;
    CCU2C _add_1_1625_add_4_8 (.A0(d_d_tmp_adj_5672[41]), .B0(d_tmp_adj_5671[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[42]), .B1(d_tmp_adj_5671[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15919), .COUT(n15920), .S0(n168_adj_5348), 
          .S1(n165_adj_5347));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_6 (.A0(d_d_tmp_adj_5672[39]), .B0(d_tmp_adj_5671[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[40]), .B1(d_tmp_adj_5671[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15918), .COUT(n15919), .S0(n174_adj_5350), 
          .S1(n171_adj_5349));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_4 (.A0(d_d_tmp_adj_5672[37]), .B0(d_tmp_adj_5671[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[38]), .B1(d_tmp_adj_5671[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15917), .COUT(n15918), .S0(n180_adj_5352), 
          .S1(n177_adj_5351));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5672[36]), .B1(d_tmp_adj_5671[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15917), .S1(n183_adj_5353));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1625_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1625_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_38 (.A0(d_d7_adj_5681[35]), .B0(d7_adj_5680[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15916), .S0(d8_71__N_1603_adj_5707[35]), 
          .S1(cout_adj_5303));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1604_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_36 (.A0(d_d7_adj_5681[33]), .B0(d7_adj_5680[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[34]), .B1(d7_adj_5680[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15915), .COUT(n15916), .S0(d8_71__N_1603_adj_5707[33]), 
          .S1(d8_71__N_1603_adj_5707[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_34 (.A0(d_d7_adj_5681[31]), .B0(d7_adj_5680[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[32]), .B1(d7_adj_5680[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15914), .COUT(n15915), .S0(d8_71__N_1603_adj_5707[31]), 
          .S1(d8_71__N_1603_adj_5707[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_32 (.A0(d_d7_adj_5681[29]), .B0(d7_adj_5680[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[30]), .B1(d7_adj_5680[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15913), .COUT(n15914), .S0(d8_71__N_1603_adj_5707[29]), 
          .S1(d8_71__N_1603_adj_5707[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_30 (.A0(d_d7_adj_5681[27]), .B0(d7_adj_5680[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[28]), .B1(d7_adj_5680[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15912), .COUT(n15913), .S0(d8_71__N_1603_adj_5707[27]), 
          .S1(d8_71__N_1603_adj_5707[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_28 (.A0(d_d7_adj_5681[25]), .B0(d7_adj_5680[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[26]), .B1(d7_adj_5680[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15911), .COUT(n15912), .S0(d8_71__N_1603_adj_5707[25]), 
          .S1(d8_71__N_1603_adj_5707[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_26 (.A0(d_d7_adj_5681[23]), .B0(d7_adj_5680[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[24]), .B1(d7_adj_5680[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15910), .COUT(n15911), .S0(d8_71__N_1603_adj_5707[23]), 
          .S1(d8_71__N_1603_adj_5707[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_24 (.A0(d_d7_adj_5681[21]), .B0(d7_adj_5680[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[22]), .B1(d7_adj_5680[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15909), .COUT(n15910), .S0(d8_71__N_1603_adj_5707[21]), 
          .S1(d8_71__N_1603_adj_5707[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_22 (.A0(d_d7_adj_5681[19]), .B0(d7_adj_5680[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[20]), .B1(d7_adj_5680[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15908), .COUT(n15909), .S0(d8_71__N_1603_adj_5707[19]), 
          .S1(d8_71__N_1603_adj_5707[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_20 (.A0(d_d7_adj_5681[17]), .B0(d7_adj_5680[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[18]), .B1(d7_adj_5680[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15907), .COUT(n15908), .S0(d8_71__N_1603_adj_5707[17]), 
          .S1(d8_71__N_1603_adj_5707[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_18 (.A0(d_d7_adj_5681[15]), .B0(d7_adj_5680[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[16]), .B1(d7_adj_5680[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15906), .COUT(n15907), .S0(d8_71__N_1603_adj_5707[15]), 
          .S1(d8_71__N_1603_adj_5707[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_16 (.A0(d_d7_adj_5681[13]), .B0(d7_adj_5680[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[14]), .B1(d7_adj_5680[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15905), .COUT(n15906), .S0(d8_71__N_1603_adj_5707[13]), 
          .S1(d8_71__N_1603_adj_5707[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_14 (.A0(d_d7_adj_5681[11]), .B0(d7_adj_5680[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[12]), .B1(d7_adj_5680[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15904), .COUT(n15905), .S0(d8_71__N_1603_adj_5707[11]), 
          .S1(d8_71__N_1603_adj_5707[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_12 (.A0(d_d7_adj_5681[9]), .B0(d7_adj_5680[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[10]), .B1(d7_adj_5680[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15903), .COUT(n15904), .S0(d8_71__N_1603_adj_5707[9]), 
          .S1(d8_71__N_1603_adj_5707[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_10 (.A0(d_d7_adj_5681[7]), .B0(d7_adj_5680[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[8]), .B1(d7_adj_5680[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15902), .COUT(n15903), .S0(d8_71__N_1603_adj_5707[7]), 
          .S1(d8_71__N_1603_adj_5707[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_8 (.A0(d_d7_adj_5681[5]), .B0(d7_adj_5680[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[6]), .B1(d7_adj_5680[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15901), .COUT(n15902), .S0(d8_71__N_1603_adj_5707[5]), 
          .S1(d8_71__N_1603_adj_5707[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_6 (.A0(d_d7_adj_5681[3]), .B0(d7_adj_5680[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[4]), .B1(d7_adj_5680[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15900), .COUT(n15901), .S0(d8_71__N_1603_adj_5707[3]), 
          .S1(d8_71__N_1603_adj_5707[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_4 (.A0(d_d7_adj_5681[1]), .B0(d7_adj_5680[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[2]), .B1(d7_adj_5680[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15899), .COUT(n15900), .S0(d8_71__N_1603_adj_5707[1]), 
          .S1(d8_71__N_1603_adj_5707[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5681[0]), .B1(d7_adj_5680[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15899), .S1(d8_71__N_1603_adj_5707[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1604_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_37 (.A0(d4[70]), .B0(cout_adj_5088), .C0(n81_adj_5449), 
          .D0(d5[70]), .A1(d4[71]), .B1(cout_adj_5088), .C1(n78_adj_5448), 
          .D1(d5[71]), .CIN(n15897), .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_35 (.A0(d4[68]), .B0(cout_adj_5088), .C0(n87_adj_5451), 
          .D0(d5[68]), .A1(d4[69]), .B1(cout_adj_5088), .C1(n84_adj_5450), 
          .D1(d5[69]), .CIN(n15896), .COUT(n15897), .S0(d5_71__N_706[68]), 
          .S1(d5_71__N_706[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_33 (.A0(d4[66]), .B0(cout_adj_5088), .C0(n93_adj_5453), 
          .D0(d5[66]), .A1(d4[67]), .B1(cout_adj_5088), .C1(n90_adj_5452), 
          .D1(d5[67]), .CIN(n15895), .COUT(n15896), .S0(d5_71__N_706[66]), 
          .S1(d5_71__N_706[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_31 (.A0(d4[64]), .B0(cout_adj_5088), .C0(n99_adj_5455), 
          .D0(d5[64]), .A1(d4[65]), .B1(cout_adj_5088), .C1(n96_adj_5454), 
          .D1(d5[65]), .CIN(n15894), .COUT(n15895), .S0(d5_71__N_706[64]), 
          .S1(d5_71__N_706[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_29 (.A0(d4[62]), .B0(cout_adj_5088), .C0(n105_adj_5457), 
          .D0(d5[62]), .A1(d4[63]), .B1(cout_adj_5088), .C1(n102_adj_5456), 
          .D1(d5[63]), .CIN(n15893), .COUT(n15894), .S0(d5_71__N_706[62]), 
          .S1(d5_71__N_706[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_27 (.A0(d4[60]), .B0(cout_adj_5088), .C0(n111_adj_5459), 
          .D0(d5[60]), .A1(d4[61]), .B1(cout_adj_5088), .C1(n108_adj_5458), 
          .D1(d5[61]), .CIN(n15892), .COUT(n15893), .S0(d5_71__N_706[60]), 
          .S1(d5_71__N_706[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_25 (.A0(d4[58]), .B0(cout_adj_5088), .C0(n117_adj_5461), 
          .D0(d5[58]), .A1(d4[59]), .B1(cout_adj_5088), .C1(n114_adj_5460), 
          .D1(d5[59]), .CIN(n15891), .COUT(n15892), .S0(d5_71__N_706[58]), 
          .S1(d5_71__N_706[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_23 (.A0(d4[56]), .B0(cout_adj_5088), .C0(n123_adj_5463), 
          .D0(d5[56]), .A1(d4[57]), .B1(cout_adj_5088), .C1(n120_adj_5462), 
          .D1(d5[57]), .CIN(n15890), .COUT(n15891), .S0(d5_71__N_706[56]), 
          .S1(d5_71__N_706[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_21 (.A0(d4[54]), .B0(cout_adj_5088), .C0(n129_adj_5465), 
          .D0(d5[54]), .A1(d4[55]), .B1(cout_adj_5088), .C1(n126_adj_5464), 
          .D1(d5[55]), .CIN(n15889), .COUT(n15890), .S0(d5_71__N_706[54]), 
          .S1(d5_71__N_706[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_19 (.A0(d4[52]), .B0(cout_adj_5088), .C0(n135_adj_5467), 
          .D0(d5[52]), .A1(d4[53]), .B1(cout_adj_5088), .C1(n132_adj_5466), 
          .D1(d5[53]), .CIN(n15888), .COUT(n15889), .S0(d5_71__N_706[52]), 
          .S1(d5_71__N_706[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_17 (.A0(d4[50]), .B0(cout_adj_5088), .C0(n141_adj_5469), 
          .D0(d5[50]), .A1(d4[51]), .B1(cout_adj_5088), .C1(n138_adj_5468), 
          .D1(d5[51]), .CIN(n15887), .COUT(n15888), .S0(d5_71__N_706[50]), 
          .S1(d5_71__N_706[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_15 (.A0(d4[48]), .B0(cout_adj_5088), .C0(n147_adj_5471), 
          .D0(d5[48]), .A1(d4[49]), .B1(cout_adj_5088), .C1(n144_adj_5470), 
          .D1(d5[49]), .CIN(n15886), .COUT(n15887), .S0(d5_71__N_706[48]), 
          .S1(d5_71__N_706[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_13 (.A0(d4[46]), .B0(cout_adj_5088), .C0(n153_adj_5473), 
          .D0(d5[46]), .A1(d4[47]), .B1(cout_adj_5088), .C1(n150_adj_5472), 
          .D1(d5[47]), .CIN(n15885), .COUT(n15886), .S0(d5_71__N_706[46]), 
          .S1(d5_71__N_706[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_11 (.A0(d4[44]), .B0(cout_adj_5088), .C0(n159_adj_5475), 
          .D0(d5[44]), .A1(d4[45]), .B1(cout_adj_5088), .C1(n156_adj_5474), 
          .D1(d5[45]), .CIN(n15884), .COUT(n15885), .S0(d5_71__N_706[44]), 
          .S1(d5_71__N_706[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_9 (.A0(d4[42]), .B0(cout_adj_5088), .C0(n165_adj_5477), 
          .D0(d5[42]), .A1(d4[43]), .B1(cout_adj_5088), .C1(n162_adj_5476), 
          .D1(d5[43]), .CIN(n15883), .COUT(n15884), .S0(d5_71__N_706[42]), 
          .S1(d5_71__N_706[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_7 (.A0(d4[40]), .B0(cout_adj_5088), .C0(n171_adj_5479), 
          .D0(d5[40]), .A1(d4[41]), .B1(cout_adj_5088), .C1(n168_adj_5478), 
          .D1(d5[41]), .CIN(n15882), .COUT(n15883), .S0(d5_71__N_706[40]), 
          .S1(d5_71__N_706[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_5 (.A0(d4[38]), .B0(cout_adj_5088), .C0(n177_adj_5481), 
          .D0(d5[38]), .A1(d4[39]), .B1(cout_adj_5088), .C1(n174_adj_5480), 
          .D1(d5[39]), .CIN(n15881), .COUT(n15882), .S0(d5_71__N_706[38]), 
          .S1(d5_71__N_706[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_3 (.A0(d4[36]), .B0(cout_adj_5088), .C0(n183_adj_5483), 
          .D0(d5[36]), .A1(d4[37]), .B1(cout_adj_5088), .C1(n180_adj_5482), 
          .D1(d5[37]), .CIN(n15880), .COUT(n15881), .S0(d5_71__N_706[36]), 
          .S1(d5_71__N_706[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5088), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15880));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1505_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1505_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_38 (.A0(d_d_tmp[35]), .B0(d_tmp[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15876), .S0(d6_71__N_1459[35]), .S1(cout_adj_5496));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1529_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_36 (.A0(d_d_tmp[33]), .B0(d_tmp[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[34]), .B1(d_tmp[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15875), .COUT(n15876), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_34 (.A0(d_d_tmp[31]), .B0(d_tmp[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[32]), .B1(d_tmp[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15874), .COUT(n15875), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_32 (.A0(d_d_tmp[29]), .B0(d_tmp[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[30]), .B1(d_tmp[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15873), .COUT(n15874), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_30 (.A0(d_d_tmp[27]), .B0(d_tmp[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[28]), .B1(d_tmp[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15872), .COUT(n15873), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_28 (.A0(d_d_tmp[25]), .B0(d_tmp[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[26]), .B1(d_tmp[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15871), .COUT(n15872), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_26 (.A0(d_d_tmp[23]), .B0(d_tmp[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[24]), .B1(d_tmp[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15870), .COUT(n15871), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_24 (.A0(d_d_tmp[21]), .B0(d_tmp[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[22]), .B1(d_tmp[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15869), .COUT(n15870), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_22 (.A0(d_d_tmp[19]), .B0(d_tmp[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[20]), .B1(d_tmp[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15868), .COUT(n15869), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_20 (.A0(d_d_tmp[17]), .B0(d_tmp[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[18]), .B1(d_tmp[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15867), .COUT(n15868), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_18 (.A0(d_d_tmp[15]), .B0(d_tmp[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[16]), .B1(d_tmp[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15866), .COUT(n15867), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_16 (.A0(d_d_tmp[13]), .B0(d_tmp[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[14]), .B1(d_tmp[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15865), .COUT(n15866), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_14 (.A0(d_d_tmp[11]), .B0(d_tmp[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[12]), .B1(d_tmp[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15864), .COUT(n15865), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_12 (.A0(d_d_tmp[9]), .B0(d_tmp[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[10]), .B1(d_tmp[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15863), .COUT(n15864), .S0(d6_71__N_1459[9]), 
          .S1(d6_71__N_1459[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_10 (.A0(d_d_tmp[7]), .B0(d_tmp[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[8]), .B1(d_tmp[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15862), .COUT(n15863), .S0(d6_71__N_1459[7]), 
          .S1(d6_71__N_1459[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_8 (.A0(d_d_tmp[5]), .B0(d_tmp[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[6]), .B1(d_tmp[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15861), .COUT(n15862), .S0(d6_71__N_1459[5]), 
          .S1(d6_71__N_1459[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_6 (.A0(d_d_tmp[3]), .B0(d_tmp[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[4]), .B1(d_tmp[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15860), .COUT(n15861), .S0(d6_71__N_1459[3]), 
          .S1(d6_71__N_1459[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_4 (.A0(d_d_tmp[1]), .B0(d_tmp[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[2]), .B1(d_tmp[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15859), .COUT(n15860), .S0(d6_71__N_1459[1]), 
          .S1(d6_71__N_1459[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1529_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[0]), .B1(d_tmp[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15859), .S1(d6_71__N_1459[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1529_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1529_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1529_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_37 (.A0(d3[70]), .B0(cout_adj_5087), .C0(n81_adj_5268), 
          .D0(d4[70]), .A1(d3[71]), .B1(cout_adj_5087), .C1(n78_adj_5267), 
          .D1(d4[71]), .CIN(n15857), .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_35 (.A0(d3[68]), .B0(cout_adj_5087), .C0(n87_adj_5270), 
          .D0(d4[68]), .A1(d3[69]), .B1(cout_adj_5087), .C1(n84_adj_5269), 
          .D1(d4[69]), .CIN(n15856), .COUT(n15857), .S0(d4_71__N_634[68]), 
          .S1(d4_71__N_634[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_33 (.A0(d3[66]), .B0(cout_adj_5087), .C0(n93_adj_5272), 
          .D0(d4[66]), .A1(d3[67]), .B1(cout_adj_5087), .C1(n90_adj_5271), 
          .D1(d4[67]), .CIN(n15855), .COUT(n15856), .S0(d4_71__N_634[66]), 
          .S1(d4_71__N_634[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_31 (.A0(d3[64]), .B0(cout_adj_5087), .C0(n99_adj_5274), 
          .D0(d4[64]), .A1(d3[65]), .B1(cout_adj_5087), .C1(n96_adj_5273), 
          .D1(d4[65]), .CIN(n15854), .COUT(n15855), .S0(d4_71__N_634[64]), 
          .S1(d4_71__N_634[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_29 (.A0(d3[62]), .B0(cout_adj_5087), .C0(n105_adj_5276), 
          .D0(d4[62]), .A1(d3[63]), .B1(cout_adj_5087), .C1(n102_adj_5275), 
          .D1(d4[63]), .CIN(n15853), .COUT(n15854), .S0(d4_71__N_634[62]), 
          .S1(d4_71__N_634[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_27 (.A0(d3[60]), .B0(cout_adj_5087), .C0(n111_adj_5278), 
          .D0(d4[60]), .A1(d3[61]), .B1(cout_adj_5087), .C1(n108_adj_5277), 
          .D1(d4[61]), .CIN(n15852), .COUT(n15853), .S0(d4_71__N_634[60]), 
          .S1(d4_71__N_634[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_25 (.A0(d3[58]), .B0(cout_adj_5087), .C0(n117_adj_5280), 
          .D0(d4[58]), .A1(d3[59]), .B1(cout_adj_5087), .C1(n114_adj_5279), 
          .D1(d4[59]), .CIN(n15851), .COUT(n15852), .S0(d4_71__N_634[58]), 
          .S1(d4_71__N_634[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_23 (.A0(d3[56]), .B0(cout_adj_5087), .C0(n123_adj_5282), 
          .D0(d4[56]), .A1(d3[57]), .B1(cout_adj_5087), .C1(n120_adj_5281), 
          .D1(d4[57]), .CIN(n15850), .COUT(n15851), .S0(d4_71__N_634[56]), 
          .S1(d4_71__N_634[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_21 (.A0(d3[54]), .B0(cout_adj_5087), .C0(n129_adj_5284), 
          .D0(d4[54]), .A1(d3[55]), .B1(cout_adj_5087), .C1(n126_adj_5283), 
          .D1(d4[55]), .CIN(n15849), .COUT(n15850), .S0(d4_71__N_634[54]), 
          .S1(d4_71__N_634[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_19 (.A0(d3[52]), .B0(cout_adj_5087), .C0(n135_adj_5286), 
          .D0(d4[52]), .A1(d3[53]), .B1(cout_adj_5087), .C1(n132_adj_5285), 
          .D1(d4[53]), .CIN(n15848), .COUT(n15849), .S0(d4_71__N_634[52]), 
          .S1(d4_71__N_634[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_17 (.A0(d3[50]), .B0(cout_adj_5087), .C0(n141_adj_5288), 
          .D0(d4[50]), .A1(d3[51]), .B1(cout_adj_5087), .C1(n138_adj_5287), 
          .D1(d4[51]), .CIN(n15847), .COUT(n15848), .S0(d4_71__N_634[50]), 
          .S1(d4_71__N_634[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_15 (.A0(d3[48]), .B0(cout_adj_5087), .C0(n147_adj_5290), 
          .D0(d4[48]), .A1(d3[49]), .B1(cout_adj_5087), .C1(n144_adj_5289), 
          .D1(d4[49]), .CIN(n15846), .COUT(n15847), .S0(d4_71__N_634[48]), 
          .S1(d4_71__N_634[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_13 (.A0(d3[46]), .B0(cout_adj_5087), .C0(n153_adj_5292), 
          .D0(d4[46]), .A1(d3[47]), .B1(cout_adj_5087), .C1(n150_adj_5291), 
          .D1(d4[47]), .CIN(n15845), .COUT(n15846), .S0(d4_71__N_634[46]), 
          .S1(d4_71__N_634[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_11 (.A0(d3[44]), .B0(cout_adj_5087), .C0(n159_adj_5294), 
          .D0(d4[44]), .A1(d3[45]), .B1(cout_adj_5087), .C1(n156_adj_5293), 
          .D1(d4[45]), .CIN(n15844), .COUT(n15845), .S0(d4_71__N_634[44]), 
          .S1(d4_71__N_634[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_9 (.A0(d3[42]), .B0(cout_adj_5087), .C0(n165_adj_5296), 
          .D0(d4[42]), .A1(d3[43]), .B1(cout_adj_5087), .C1(n162_adj_5295), 
          .D1(d4[43]), .CIN(n15843), .COUT(n15844), .S0(d4_71__N_634[42]), 
          .S1(d4_71__N_634[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_7 (.A0(d3[40]), .B0(cout_adj_5087), .C0(n171_adj_5298), 
          .D0(d4[40]), .A1(d3[41]), .B1(cout_adj_5087), .C1(n168_adj_5297), 
          .D1(d4[41]), .CIN(n15842), .COUT(n15843), .S0(d4_71__N_634[40]), 
          .S1(d4_71__N_634[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_5 (.A0(d3[38]), .B0(cout_adj_5087), .C0(n177_adj_5300), 
          .D0(d4[38]), .A1(d3[39]), .B1(cout_adj_5087), .C1(n174_adj_5299), 
          .D1(d4[39]), .CIN(n15841), .COUT(n15842), .S0(d4_71__N_634[38]), 
          .S1(d4_71__N_634[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_3 (.A0(d3[36]), .B0(cout_adj_5087), .C0(n183_adj_5302), 
          .D0(d4[36]), .A1(d3[37]), .B1(cout_adj_5087), .C1(n180_adj_5301), 
          .D1(d4[37]), .CIN(n15840), .COUT(n15841), .S0(d4_71__N_634[36]), 
          .S1(d4_71__N_634[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5087), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15840));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1508_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1508_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_37 (.A0(d2[70]), .B0(cout_adj_4736), .C0(n81_adj_5232), 
          .D0(d3[70]), .A1(d2[71]), .B1(cout_adj_4736), .C1(n78_adj_5231), 
          .D1(d3[71]), .CIN(n15835), .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_35 (.A0(d2[68]), .B0(cout_adj_4736), .C0(n87_adj_5234), 
          .D0(d3[68]), .A1(d2[69]), .B1(cout_adj_4736), .C1(n84_adj_5233), 
          .D1(d3[69]), .CIN(n15834), .COUT(n15835), .S0(d3_71__N_562[68]), 
          .S1(d3_71__N_562[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_33 (.A0(d2[66]), .B0(cout_adj_4736), .C0(n93_adj_5236), 
          .D0(d3[66]), .A1(d2[67]), .B1(cout_adj_4736), .C1(n90_adj_5235), 
          .D1(d3[67]), .CIN(n15833), .COUT(n15834), .S0(d3_71__N_562[66]), 
          .S1(d3_71__N_562[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_31 (.A0(d2[64]), .B0(cout_adj_4736), .C0(n99_adj_5238), 
          .D0(d3[64]), .A1(d2[65]), .B1(cout_adj_4736), .C1(n96_adj_5237), 
          .D1(d3[65]), .CIN(n15832), .COUT(n15833), .S0(d3_71__N_562[64]), 
          .S1(d3_71__N_562[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_29 (.A0(d2[62]), .B0(cout_adj_4736), .C0(n105_adj_5240), 
          .D0(d3[62]), .A1(d2[63]), .B1(cout_adj_4736), .C1(n102_adj_5239), 
          .D1(d3[63]), .CIN(n15831), .COUT(n15832), .S0(d3_71__N_562[62]), 
          .S1(d3_71__N_562[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_27 (.A0(d2[60]), .B0(cout_adj_4736), .C0(n111_adj_5242), 
          .D0(d3[60]), .A1(d2[61]), .B1(cout_adj_4736), .C1(n108_adj_5241), 
          .D1(d3[61]), .CIN(n15830), .COUT(n15831), .S0(d3_71__N_562[60]), 
          .S1(d3_71__N_562[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_25 (.A0(d2[58]), .B0(cout_adj_4736), .C0(n117_adj_5244), 
          .D0(d3[58]), .A1(d2[59]), .B1(cout_adj_4736), .C1(n114_adj_5243), 
          .D1(d3[59]), .CIN(n15829), .COUT(n15830), .S0(d3_71__N_562[58]), 
          .S1(d3_71__N_562[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_23 (.A0(d2[56]), .B0(cout_adj_4736), .C0(n123_adj_5246), 
          .D0(d3[56]), .A1(d2[57]), .B1(cout_adj_4736), .C1(n120_adj_5245), 
          .D1(d3[57]), .CIN(n15828), .COUT(n15829), .S0(d3_71__N_562[56]), 
          .S1(d3_71__N_562[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_21 (.A0(d2[54]), .B0(cout_adj_4736), .C0(n129_adj_5248), 
          .D0(d3[54]), .A1(d2[55]), .B1(cout_adj_4736), .C1(n126_adj_5247), 
          .D1(d3[55]), .CIN(n15827), .COUT(n15828), .S0(d3_71__N_562[54]), 
          .S1(d3_71__N_562[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_19 (.A0(d2[52]), .B0(cout_adj_4736), .C0(n135_adj_5250), 
          .D0(d3[52]), .A1(d2[53]), .B1(cout_adj_4736), .C1(n132_adj_5249), 
          .D1(d3[53]), .CIN(n15826), .COUT(n15827), .S0(d3_71__N_562[52]), 
          .S1(d3_71__N_562[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_17 (.A0(d2[50]), .B0(cout_adj_4736), .C0(n141_adj_5252), 
          .D0(d3[50]), .A1(d2[51]), .B1(cout_adj_4736), .C1(n138_adj_5251), 
          .D1(d3[51]), .CIN(n15825), .COUT(n15826), .S0(d3_71__N_562[50]), 
          .S1(d3_71__N_562[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_15 (.A0(d2[48]), .B0(cout_adj_4736), .C0(n147_adj_5254), 
          .D0(d3[48]), .A1(d2[49]), .B1(cout_adj_4736), .C1(n144_adj_5253), 
          .D1(d3[49]), .CIN(n15824), .COUT(n15825), .S0(d3_71__N_562[48]), 
          .S1(d3_71__N_562[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_13 (.A0(d2[46]), .B0(cout_adj_4736), .C0(n153_adj_5256), 
          .D0(d3[46]), .A1(d2[47]), .B1(cout_adj_4736), .C1(n150_adj_5255), 
          .D1(d3[47]), .CIN(n15823), .COUT(n15824), .S0(d3_71__N_562[46]), 
          .S1(d3_71__N_562[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_11 (.A0(d2[44]), .B0(cout_adj_4736), .C0(n159_adj_5258), 
          .D0(d3[44]), .A1(d2[45]), .B1(cout_adj_4736), .C1(n156_adj_5257), 
          .D1(d3[45]), .CIN(n15822), .COUT(n15823), .S0(d3_71__N_562[44]), 
          .S1(d3_71__N_562[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_9 (.A0(d2[42]), .B0(cout_adj_4736), .C0(n165_adj_5260), 
          .D0(d3[42]), .A1(d2[43]), .B1(cout_adj_4736), .C1(n162_adj_5259), 
          .D1(d3[43]), .CIN(n15821), .COUT(n15822), .S0(d3_71__N_562[42]), 
          .S1(d3_71__N_562[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_7 (.A0(d2[40]), .B0(cout_adj_4736), .C0(n171_adj_5262), 
          .D0(d3[40]), .A1(d2[41]), .B1(cout_adj_4736), .C1(n168_adj_5261), 
          .D1(d3[41]), .CIN(n15820), .COUT(n15821), .S0(d3_71__N_562[40]), 
          .S1(d3_71__N_562[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_5 (.A0(d2[38]), .B0(cout_adj_4736), .C0(n177_adj_5264), 
          .D0(d3[38]), .A1(d2[39]), .B1(cout_adj_4736), .C1(n174_adj_5263), 
          .D1(d3[39]), .CIN(n15819), .COUT(n15820), .S0(d3_71__N_562[38]), 
          .S1(d3_71__N_562[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_3 (.A0(d2[36]), .B0(cout_adj_4736), .C0(n183_adj_5266), 
          .D0(d3[36]), .A1(d2[37]), .B1(cout_adj_4736), .C1(n180_adj_5265), 
          .D1(d3[37]), .CIN(n15818), .COUT(n15819), .S0(d3_71__N_562[36]), 
          .S1(d3_71__N_562[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4736), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15818));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1511_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1511_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_38 (.A0(d2[71]), .B0(d1[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15814), .S0(n78_adj_5193));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1556_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_36 (.A0(d2[69]), .B0(d1[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[70]), .B1(d1[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15813), .COUT(n15814), .S0(n84_adj_5195), .S1(n81_adj_5194));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_34 (.A0(d2[67]), .B0(d1[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[68]), .B1(d1[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15812), .COUT(n15813), .S0(n90_adj_5197), .S1(n87_adj_5196));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_32 (.A0(d2[65]), .B0(d1[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[66]), .B1(d1[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15811), .COUT(n15812), .S0(n96_adj_5199), .S1(n93_adj_5198));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_30 (.A0(d2[63]), .B0(d1[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[64]), .B1(d1[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15810), .COUT(n15811), .S0(n102_adj_5201), .S1(n99_adj_5200));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_28 (.A0(d2[61]), .B0(d1[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[62]), .B1(d1[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15809), .COUT(n15810), .S0(n108_adj_5203), .S1(n105_adj_5202));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_26 (.A0(d2[59]), .B0(d1[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[60]), .B1(d1[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15808), .COUT(n15809), .S0(n114_adj_5205), .S1(n111_adj_5204));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_24 (.A0(d2[57]), .B0(d1[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[58]), .B1(d1[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15807), .COUT(n15808), .S0(n120_adj_5207), .S1(n117_adj_5206));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_22 (.A0(d2[55]), .B0(d1[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[56]), .B1(d1[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15806), .COUT(n15807), .S0(n126_adj_5209), .S1(n123_adj_5208));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_20 (.A0(d2[53]), .B0(d1[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[54]), .B1(d1[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15805), .COUT(n15806), .S0(n132_adj_5211), .S1(n129_adj_5210));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_18 (.A0(d2[51]), .B0(d1[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[52]), .B1(d1[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15804), .COUT(n15805), .S0(n138_adj_5213), .S1(n135_adj_5212));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_16 (.A0(d2[49]), .B0(d1[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[50]), .B1(d1[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15803), .COUT(n15804), .S0(n144_adj_5215), .S1(n141_adj_5214));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_14 (.A0(d2[47]), .B0(d1[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[48]), .B1(d1[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15802), .COUT(n15803), .S0(n150_adj_5217), .S1(n147_adj_5216));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_12 (.A0(d2[45]), .B0(d1[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[46]), .B1(d1[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15801), .COUT(n15802), .S0(n156_adj_5219), .S1(n153_adj_5218));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_10 (.A0(d2[43]), .B0(d1[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[44]), .B1(d1[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15800), .COUT(n15801), .S0(n162_adj_5221), .S1(n159_adj_5220));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_8 (.A0(d2[41]), .B0(d1[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[42]), .B1(d1[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15799), .COUT(n15800), .S0(n168_adj_5223), .S1(n165_adj_5222));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_6 (.A0(d2[39]), .B0(d1[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[40]), .B1(d1[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15798), .COUT(n15799), .S0(n174_adj_5225), .S1(n171_adj_5224));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_4 (.A0(d2[37]), .B0(d1[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[38]), .B1(d1[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15797), .COUT(n15798), .S0(n180_adj_5227), .S1(n177_adj_5226));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[36]), .B1(d1[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15797), .S1(n183_adj_5228));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1556_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1556_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_38 (.A0(d_d9_adj_5685[35]), .B0(d9_adj_5684[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15796), .S1(cout_adj_5229));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1598_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_36 (.A0(d_d9_adj_5685[33]), .B0(d9_adj_5684[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[34]), .B1(d9_adj_5684[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15795), .COUT(n15796));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_34 (.A0(d_d9_adj_5685[31]), .B0(d9_adj_5684[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[32]), .B1(d9_adj_5684[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15794), .COUT(n15795));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_32 (.A0(d_d9_adj_5685[29]), .B0(d9_adj_5684[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[30]), .B1(d9_adj_5684[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15793), .COUT(n15794));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_30 (.A0(d_d9_adj_5685[27]), .B0(d9_adj_5684[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[28]), .B1(d9_adj_5684[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15792), .COUT(n15793));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_28 (.A0(d_d9_adj_5685[25]), .B0(d9_adj_5684[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[26]), .B1(d9_adj_5684[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15791), .COUT(n15792));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_26 (.A0(d_d9_adj_5685[23]), .B0(d9_adj_5684[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[24]), .B1(d9_adj_5684[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15790), .COUT(n15791));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_24 (.A0(d_d9_adj_5685[21]), .B0(d9_adj_5684[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[22]), .B1(d9_adj_5684[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15789), .COUT(n15790));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_22 (.A0(d_d9_adj_5685[19]), .B0(d9_adj_5684[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[20]), .B1(d9_adj_5684[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15788), .COUT(n15789));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_20 (.A0(d_d9_adj_5685[17]), .B0(d9_adj_5684[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[18]), .B1(d9_adj_5684[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15787), .COUT(n15788));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_18 (.A0(d_d9_adj_5685[15]), .B0(d9_adj_5684[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[16]), .B1(d9_adj_5684[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15786), .COUT(n15787));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_16 (.A0(d_d9_adj_5685[13]), .B0(d9_adj_5684[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[14]), .B1(d9_adj_5684[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15785), .COUT(n15786));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_14 (.A0(d_d9_adj_5685[11]), .B0(d9_adj_5684[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[12]), .B1(d9_adj_5684[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15784), .COUT(n15785));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_12 (.A0(d_d9_adj_5685[9]), .B0(d9_adj_5684[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[10]), .B1(d9_adj_5684[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15783), .COUT(n15784));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_10 (.A0(d_d9_adj_5685[7]), .B0(d9_adj_5684[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[8]), .B1(d9_adj_5684[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15782), .COUT(n15783));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_8 (.A0(d_d9_adj_5685[5]), .B0(d9_adj_5684[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[6]), .B1(d9_adj_5684[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15781), .COUT(n15782));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_8.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i2 (.D(n123_adj_5190), .CK(CIC1_out_clkSin), .Q(ISquare[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i2.GSR = "ENABLED";
    LUT4 i5662_2_lut (.A(phase_inc_carrGen1[0]), .B(phase_accum_adj_5665[0]), 
         .Z(n321)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5662_2_lut.init = 16'h6666;
    LUT4 i2490_4_lut (.A(n133_adj_5391), .B(n127), .C(led_c_3), .D(n18141), 
         .Z(n12221)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2490_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n18138), .B(n18267), .C(n235), .D(led_c_3), 
         .Z(n11999)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_3_lut_3_lut_4_lut.init = 16'hf088;
    LUT4 i5619_2_lut (.A(d1[0]), .B(MixerOutSin[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5619_2_lut.init = 16'h6666;
    CCU2C _add_1_1598_add_4_6 (.A0(d_d9_adj_5685[3]), .B0(d9_adj_5684[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[4]), .B1(d9_adj_5684[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15780), .COUT(n15781));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_4 (.A0(d_d9_adj_5685[1]), .B0(d9_adj_5684[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[2]), .B1(d9_adj_5684[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15779), .COUT(n15780));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1598_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1598_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5685[0]), .B1(d9_adj_5684[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15779));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1598_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1598_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1598_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1598_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_38 (.A0(d_d8_adj_5683[35]), .B0(d8_adj_5682[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15778), .S0(d9_71__N_1675_adj_5708[35]), 
          .S1(cout_adj_5230));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1601_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_36 (.A0(d_d8_adj_5683[33]), .B0(d8_adj_5682[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[34]), .B1(d8_adj_5682[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15777), .COUT(n15778), .S0(d9_71__N_1675_adj_5708[33]), 
          .S1(d9_71__N_1675_adj_5708[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_34 (.A0(d_d8_adj_5683[31]), .B0(d8_adj_5682[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[32]), .B1(d8_adj_5682[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15776), .COUT(n15777), .S0(d9_71__N_1675_adj_5708[31]), 
          .S1(d9_71__N_1675_adj_5708[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_32 (.A0(d_d8_adj_5683[29]), .B0(d8_adj_5682[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[30]), .B1(d8_adj_5682[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15775), .COUT(n15776), .S0(d9_71__N_1675_adj_5708[29]), 
          .S1(d9_71__N_1675_adj_5708[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_30 (.A0(d_d8_adj_5683[27]), .B0(d8_adj_5682[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[28]), .B1(d8_adj_5682[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15774), .COUT(n15775), .S0(d9_71__N_1675_adj_5708[27]), 
          .S1(d9_71__N_1675_adj_5708[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_28 (.A0(d_d8_adj_5683[25]), .B0(d8_adj_5682[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[26]), .B1(d8_adj_5682[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15773), .COUT(n15774), .S0(d9_71__N_1675_adj_5708[25]), 
          .S1(d9_71__N_1675_adj_5708[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_26 (.A0(d_d8_adj_5683[23]), .B0(d8_adj_5682[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[24]), .B1(d8_adj_5682[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15772), .COUT(n15773), .S0(d9_71__N_1675_adj_5708[23]), 
          .S1(d9_71__N_1675_adj_5708[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_24 (.A0(d_d8_adj_5683[21]), .B0(d8_adj_5682[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[22]), .B1(d8_adj_5682[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15771), .COUT(n15772), .S0(d9_71__N_1675_adj_5708[21]), 
          .S1(d9_71__N_1675_adj_5708[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_22 (.A0(d_d8_adj_5683[19]), .B0(d8_adj_5682[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[20]), .B1(d8_adj_5682[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15770), .COUT(n15771), .S0(d9_71__N_1675_adj_5708[19]), 
          .S1(d9_71__N_1675_adj_5708[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_20 (.A0(d_d8_adj_5683[17]), .B0(d8_adj_5682[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[18]), .B1(d8_adj_5682[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15769), .COUT(n15770), .S0(d9_71__N_1675_adj_5708[17]), 
          .S1(d9_71__N_1675_adj_5708[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_18 (.A0(d_d8_adj_5683[15]), .B0(d8_adj_5682[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[16]), .B1(d8_adj_5682[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15768), .COUT(n15769), .S0(d9_71__N_1675_adj_5708[15]), 
          .S1(d9_71__N_1675_adj_5708[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_16 (.A0(d_d8_adj_5683[13]), .B0(d8_adj_5682[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[14]), .B1(d8_adj_5682[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15767), .COUT(n15768), .S0(d9_71__N_1675_adj_5708[13]), 
          .S1(d9_71__N_1675_adj_5708[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_14 (.A0(d_d8_adj_5683[11]), .B0(d8_adj_5682[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[12]), .B1(d8_adj_5682[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15766), .COUT(n15767), .S0(d9_71__N_1675_adj_5708[11]), 
          .S1(d9_71__N_1675_adj_5708[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_12 (.A0(d_d8_adj_5683[9]), .B0(d8_adj_5682[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[10]), .B1(d8_adj_5682[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15765), .COUT(n15766), .S0(d9_71__N_1675_adj_5708[9]), 
          .S1(d9_71__N_1675_adj_5708[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_10 (.A0(d_d8_adj_5683[7]), .B0(d8_adj_5682[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[8]), .B1(d8_adj_5682[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15764), .COUT(n15765), .S0(d9_71__N_1675_adj_5708[7]), 
          .S1(d9_71__N_1675_adj_5708[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_8 (.A0(d_d8_adj_5683[5]), .B0(d8_adj_5682[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[6]), .B1(d8_adj_5682[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15763), .COUT(n15764), .S0(d9_71__N_1675_adj_5708[5]), 
          .S1(d9_71__N_1675_adj_5708[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_6 (.A0(d_d8_adj_5683[3]), .B0(d8_adj_5682[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[4]), .B1(d8_adj_5682[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15762), .COUT(n15763), .S0(d9_71__N_1675_adj_5708[3]), 
          .S1(d9_71__N_1675_adj_5708[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_4 (.A0(d_d8_adj_5683[1]), .B0(d8_adj_5682[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[2]), .B1(d8_adj_5682[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15761), .COUT(n15762), .S0(d9_71__N_1675_adj_5708[1]), 
          .S1(d9_71__N_1675_adj_5708[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5683[0]), .B1(d8_adj_5682[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15761), .S1(d9_71__N_1675_adj_5708[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1601_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_37 (.A0(d1[70]), .B0(cout), .C0(n81_adj_5194), 
          .D0(d2[70]), .A1(d1[71]), .B1(cout), .C1(n78_adj_5193), .D1(d2[71]), 
          .CIN(n15759), .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_35 (.A0(d1[68]), .B0(cout), .C0(n87_adj_5196), 
          .D0(d2[68]), .A1(d1[69]), .B1(cout), .C1(n84_adj_5195), .D1(d2[69]), 
          .CIN(n15758), .COUT(n15759), .S0(d2_71__N_490[68]), .S1(d2_71__N_490[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_33 (.A0(d1[66]), .B0(cout), .C0(n93_adj_5198), 
          .D0(d2[66]), .A1(d1[67]), .B1(cout), .C1(n90_adj_5197), .D1(d2[67]), 
          .CIN(n15757), .COUT(n15758), .S0(d2_71__N_490[66]), .S1(d2_71__N_490[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_31 (.A0(d1[64]), .B0(cout), .C0(n99_adj_5200), 
          .D0(d2[64]), .A1(d1[65]), .B1(cout), .C1(n96_adj_5199), .D1(d2[65]), 
          .CIN(n15756), .COUT(n15757), .S0(d2_71__N_490[64]), .S1(d2_71__N_490[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_29 (.A0(d1[62]), .B0(cout), .C0(n105_adj_5202), 
          .D0(d2[62]), .A1(d1[63]), .B1(cout), .C1(n102_adj_5201), .D1(d2[63]), 
          .CIN(n15755), .COUT(n15756), .S0(d2_71__N_490[62]), .S1(d2_71__N_490[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_27 (.A0(d1[60]), .B0(cout), .C0(n111_adj_5204), 
          .D0(d2[60]), .A1(d1[61]), .B1(cout), .C1(n108_adj_5203), .D1(d2[61]), 
          .CIN(n15754), .COUT(n15755), .S0(d2_71__N_490[60]), .S1(d2_71__N_490[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_25 (.A0(d1[58]), .B0(cout), .C0(n117_adj_5206), 
          .D0(d2[58]), .A1(d1[59]), .B1(cout), .C1(n114_adj_5205), .D1(d2[59]), 
          .CIN(n15753), .COUT(n15754), .S0(d2_71__N_490[58]), .S1(d2_71__N_490[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_23 (.A0(d1[56]), .B0(cout), .C0(n123_adj_5208), 
          .D0(d2[56]), .A1(d1[57]), .B1(cout), .C1(n120_adj_5207), .D1(d2[57]), 
          .CIN(n15752), .COUT(n15753), .S0(d2_71__N_490[56]), .S1(d2_71__N_490[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_21 (.A0(d1[54]), .B0(cout), .C0(n129_adj_5210), 
          .D0(d2[54]), .A1(d1[55]), .B1(cout), .C1(n126_adj_5209), .D1(d2[55]), 
          .CIN(n15751), .COUT(n15752), .S0(d2_71__N_490[54]), .S1(d2_71__N_490[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_19 (.A0(d1[52]), .B0(cout), .C0(n135_adj_5212), 
          .D0(d2[52]), .A1(d1[53]), .B1(cout), .C1(n132_adj_5211), .D1(d2[53]), 
          .CIN(n15750), .COUT(n15751), .S0(d2_71__N_490[52]), .S1(d2_71__N_490[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_17 (.A0(d1[50]), .B0(cout), .C0(n141_adj_5214), 
          .D0(d2[50]), .A1(d1[51]), .B1(cout), .C1(n138_adj_5213), .D1(d2[51]), 
          .CIN(n15749), .COUT(n15750), .S0(d2_71__N_490[50]), .S1(d2_71__N_490[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_15 (.A0(d1[48]), .B0(cout), .C0(n147_adj_5216), 
          .D0(d2[48]), .A1(d1[49]), .B1(cout), .C1(n144_adj_5215), .D1(d2[49]), 
          .CIN(n15748), .COUT(n15749), .S0(d2_71__N_490[48]), .S1(d2_71__N_490[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_13 (.A0(d1[46]), .B0(cout), .C0(n153_adj_5218), 
          .D0(d2[46]), .A1(d1[47]), .B1(cout), .C1(n150_adj_5217), .D1(d2[47]), 
          .CIN(n15747), .COUT(n15748), .S0(d2_71__N_490[46]), .S1(d2_71__N_490[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_11 (.A0(d1[44]), .B0(cout), .C0(n159_adj_5220), 
          .D0(d2[44]), .A1(d1[45]), .B1(cout), .C1(n156_adj_5219), .D1(d2[45]), 
          .CIN(n15746), .COUT(n15747), .S0(d2_71__N_490[44]), .S1(d2_71__N_490[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_9 (.A0(d1[42]), .B0(cout), .C0(n165_adj_5222), 
          .D0(d2[42]), .A1(d1[43]), .B1(cout), .C1(n162_adj_5221), .D1(d2[43]), 
          .CIN(n15745), .COUT(n15746), .S0(d2_71__N_490[42]), .S1(d2_71__N_490[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_7 (.A0(d1[40]), .B0(cout), .C0(n171_adj_5224), 
          .D0(d2[40]), .A1(d1[41]), .B1(cout), .C1(n168_adj_5223), .D1(d2[41]), 
          .CIN(n15744), .COUT(n15745), .S0(d2_71__N_490[40]), .S1(d2_71__N_490[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_5 (.A0(d1[38]), .B0(cout), .C0(n177_adj_5226), 
          .D0(d2[38]), .A1(d1[39]), .B1(cout), .C1(n174_adj_5225), .D1(d2[39]), 
          .CIN(n15743), .COUT(n15744), .S0(d2_71__N_490[38]), .S1(d2_71__N_490[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_3 (.A0(d1[36]), .B0(cout), .C0(n183_adj_5228), 
          .D0(d2[36]), .A1(d1[37]), .B1(cout), .C1(n180_adj_5227), .D1(d2[37]), 
          .CIN(n15742), .COUT(n15743), .S0(d2_71__N_490[36]), .S1(d2_71__N_490[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1514_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1514_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1514_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15742));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1514_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1514_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1514_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1514_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_38 (.A0(d_d7_adj_5681[71]), .B0(d7_adj_5680[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15738), .S0(n78_adj_2770));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1631_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_36 (.A0(d_d7_adj_5681[69]), .B0(d7_adj_5680[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[70]), .B1(d7_adj_5680[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15737), .COUT(n15738), .S0(n84_adj_2768), 
          .S1(n81_adj_2769));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_34 (.A0(d_d7_adj_5681[67]), .B0(d7_adj_5680[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[68]), .B1(d7_adj_5680[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15736), .COUT(n15737), .S0(n90_adj_2766), 
          .S1(n87_adj_2767));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_32 (.A0(d_d7_adj_5681[65]), .B0(d7_adj_5680[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[66]), .B1(d7_adj_5680[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15735), .COUT(n15736), .S0(n96_adj_2764), 
          .S1(n93_adj_2765));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_30 (.A0(d_d7_adj_5681[63]), .B0(d7_adj_5680[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[64]), .B1(d7_adj_5680[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15734), .COUT(n15735), .S0(n102_adj_2762), 
          .S1(n99_adj_2763));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_28 (.A0(d_d7_adj_5681[61]), .B0(d7_adj_5680[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[62]), .B1(d7_adj_5680[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15733), .COUT(n15734), .S0(n108), 
          .S1(n105));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_26 (.A0(d_d7_adj_5681[59]), .B0(d7_adj_5680[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[60]), .B1(d7_adj_5680[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15732), .COUT(n15733), .S0(n114), 
          .S1(n111));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_24 (.A0(d_d7_adj_5681[57]), .B0(d7_adj_5680[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[58]), .B1(d7_adj_5680[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15731), .COUT(n15732), .S0(n120), 
          .S1(n117));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_22 (.A0(d_d7_adj_5681[55]), .B0(d7_adj_5680[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[56]), .B1(d7_adj_5680[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15730), .COUT(n15731), .S0(n126), 
          .S1(n123));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_20 (.A0(d_d7_adj_5681[53]), .B0(d7_adj_5680[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[54]), .B1(d7_adj_5680[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15729), .COUT(n15730), .S0(n132), 
          .S1(n129));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_18 (.A0(d_d7_adj_5681[51]), .B0(d7_adj_5680[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[52]), .B1(d7_adj_5680[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15728), .COUT(n15729), .S0(n138), 
          .S1(n135));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_16 (.A0(d_d7_adj_5681[49]), .B0(d7_adj_5680[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[50]), .B1(d7_adj_5680[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15727), .COUT(n15728), .S0(n144), 
          .S1(n141));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_14 (.A0(d_d7_adj_5681[47]), .B0(d7_adj_5680[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[48]), .B1(d7_adj_5680[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15726), .COUT(n15727), .S0(n150), 
          .S1(n147));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_12 (.A0(d_d7_adj_5681[45]), .B0(d7_adj_5680[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[46]), .B1(d7_adj_5680[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15725), .COUT(n15726), .S0(n156), 
          .S1(n153));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_10 (.A0(d_d7_adj_5681[43]), .B0(d7_adj_5680[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[44]), .B1(d7_adj_5680[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15724), .COUT(n15725), .S0(n162), 
          .S1(n159));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_8 (.A0(d_d7_adj_5681[41]), .B0(d7_adj_5680[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[42]), .B1(d7_adj_5680[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15723), .COUT(n15724), .S0(n168), 
          .S1(n165));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_6 (.A0(d_d7_adj_5681[39]), .B0(d7_adj_5680[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[40]), .B1(d7_adj_5680[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15722), .COUT(n15723), .S0(n174), 
          .S1(n171));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_4 (.A0(d_d7_adj_5681[37]), .B0(d7_adj_5680[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5681[38]), .B1(d7_adj_5680[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15721), .COUT(n15722), .S0(n180), 
          .S1(n177));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5681[36]), .B1(d7_adj_5680[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15721), .S1(n183));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1631_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1631_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_38 (.A0(d3[71]), .B0(d2[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15720), .S0(n78_adj_5231));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1559_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_36 (.A0(d3[69]), .B0(d2[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[70]), .B1(d2[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15719), .COUT(n15720), .S0(n84_adj_5233), .S1(n81_adj_5232));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_34 (.A0(d3[67]), .B0(d2[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[68]), .B1(d2[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15718), .COUT(n15719), .S0(n90_adj_5235), .S1(n87_adj_5234));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_32 (.A0(d3[65]), .B0(d2[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[66]), .B1(d2[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15717), .COUT(n15718), .S0(n96_adj_5237), .S1(n93_adj_5236));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_30 (.A0(d3[63]), .B0(d2[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[64]), .B1(d2[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15716), .COUT(n15717), .S0(n102_adj_5239), .S1(n99_adj_5238));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_28 (.A0(d3[61]), .B0(d2[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[62]), .B1(d2[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15715), .COUT(n15716), .S0(n108_adj_5241), .S1(n105_adj_5240));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_26 (.A0(d3[59]), .B0(d2[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[60]), .B1(d2[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15714), .COUT(n15715), .S0(n114_adj_5243), .S1(n111_adj_5242));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_24 (.A0(d3[57]), .B0(d2[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[58]), .B1(d2[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15713), .COUT(n15714), .S0(n120_adj_5245), .S1(n117_adj_5244));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_22 (.A0(d3[55]), .B0(d2[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[56]), .B1(d2[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15712), .COUT(n15713), .S0(n126_adj_5247), .S1(n123_adj_5246));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_20 (.A0(d3[53]), .B0(d2[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[54]), .B1(d2[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15711), .COUT(n15712), .S0(n132_adj_5249), .S1(n129_adj_5248));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_18 (.A0(d3[51]), .B0(d2[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[52]), .B1(d2[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15710), .COUT(n15711), .S0(n138_adj_5251), .S1(n135_adj_5250));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_16 (.A0(d3[49]), .B0(d2[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[50]), .B1(d2[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15709), .COUT(n15710), .S0(n144_adj_5253), .S1(n141_adj_5252));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_14 (.A0(d3[47]), .B0(d2[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[48]), .B1(d2[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15708), .COUT(n15709), .S0(n150_adj_5255), .S1(n147_adj_5254));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_12 (.A0(d3[45]), .B0(d2[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[46]), .B1(d2[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15707), .COUT(n15708), .S0(n156_adj_5257), .S1(n153_adj_5256));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_10 (.A0(d3[43]), .B0(d2[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[44]), .B1(d2[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15706), .COUT(n15707), .S0(n162_adj_5259), .S1(n159_adj_5258));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_8 (.A0(d3[41]), .B0(d2[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[42]), .B1(d2[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15705), .COUT(n15706), .S0(n168_adj_5261), .S1(n165_adj_5260));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_6 (.A0(d3[39]), .B0(d2[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[40]), .B1(d2[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15704), .COUT(n15705), .S0(n174_adj_5263), .S1(n171_adj_5262));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_4 (.A0(d3[37]), .B0(d2[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[38]), .B1(d2[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15703), .COUT(n15704), .S0(n180_adj_5265), .S1(n177_adj_5264));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[36]), .B1(d2[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15703), .S1(n183_adj_5266));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1559_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1559_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_37 (.A0(d7_adj_5680[70]), .B0(cout_adj_5303), 
          .C0(n81_adj_2769), .D0(n3_adj_4653), .A1(d7_adj_5680[71]), .B1(cout_adj_5303), 
          .C1(n78_adj_2770), .D1(n2_adj_4654), .CIN(n15701), .S0(d8_71__N_1603_adj_5707[70]), 
          .S1(d8_71__N_1603_adj_5707[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_35 (.A0(d7_adj_5680[68]), .B0(cout_adj_5303), 
          .C0(n87_adj_2767), .D0(n5_adj_4651), .A1(d7_adj_5680[69]), .B1(cout_adj_5303), 
          .C1(n84_adj_2768), .D1(n4_adj_4652), .CIN(n15700), .COUT(n15701), 
          .S0(d8_71__N_1603_adj_5707[68]), .S1(d8_71__N_1603_adj_5707[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_33 (.A0(d7_adj_5680[66]), .B0(cout_adj_5303), 
          .C0(n93_adj_2765), .D0(n7_adj_4649), .A1(d7_adj_5680[67]), .B1(cout_adj_5303), 
          .C1(n90_adj_2766), .D1(n6_adj_4650), .CIN(n15699), .COUT(n15700), 
          .S0(d8_71__N_1603_adj_5707[66]), .S1(d8_71__N_1603_adj_5707[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_31 (.A0(d7_adj_5680[64]), .B0(cout_adj_5303), 
          .C0(n99_adj_2763), .D0(n9_adj_4647), .A1(d7_adj_5680[65]), .B1(cout_adj_5303), 
          .C1(n96_adj_2764), .D1(n8_adj_4648), .CIN(n15698), .COUT(n15699), 
          .S0(d8_71__N_1603_adj_5707[64]), .S1(d8_71__N_1603_adj_5707[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_29 (.A0(d7_adj_5680[62]), .B0(cout_adj_5303), 
          .C0(n105), .D0(n11_adj_4645), .A1(d7_adj_5680[63]), .B1(cout_adj_5303), 
          .C1(n102_adj_2762), .D1(n10_adj_4646), .CIN(n15697), .COUT(n15698), 
          .S0(d8_71__N_1603_adj_5707[62]), .S1(d8_71__N_1603_adj_5707[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_27 (.A0(d7_adj_5680[60]), .B0(cout_adj_5303), 
          .C0(n111), .D0(n13_adj_4643), .A1(d7_adj_5680[61]), .B1(cout_adj_5303), 
          .C1(n108), .D1(n12_adj_4644), .CIN(n15696), .COUT(n15697), 
          .S0(d8_71__N_1603_adj_5707[60]), .S1(d8_71__N_1603_adj_5707[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_25 (.A0(d7_adj_5680[58]), .B0(cout_adj_5303), 
          .C0(n117), .D0(n15_adj_4641), .A1(d7_adj_5680[59]), .B1(cout_adj_5303), 
          .C1(n114), .D1(n14_adj_4642), .CIN(n15695), .COUT(n15696), 
          .S0(d8_71__N_1603_adj_5707[58]), .S1(d8_71__N_1603_adj_5707[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_23 (.A0(d7_adj_5680[56]), .B0(cout_adj_5303), 
          .C0(n123), .D0(n17_adj_4639), .A1(d7_adj_5680[57]), .B1(cout_adj_5303), 
          .C1(n120), .D1(n16_adj_4640), .CIN(n15694), .COUT(n15695), 
          .S0(d8_71__N_1603_adj_5707[56]), .S1(d8_71__N_1603_adj_5707[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_21 (.A0(d7_adj_5680[54]), .B0(cout_adj_5303), 
          .C0(n129), .D0(n19_adj_4637), .A1(d7_adj_5680[55]), .B1(cout_adj_5303), 
          .C1(n126), .D1(n18_adj_4638), .CIN(n15693), .COUT(n15694), 
          .S0(d8_71__N_1603_adj_5707[54]), .S1(d8_71__N_1603_adj_5707[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_19 (.A0(d7_adj_5680[52]), .B0(cout_adj_5303), 
          .C0(n135), .D0(n21_adj_4635), .A1(d7_adj_5680[53]), .B1(cout_adj_5303), 
          .C1(n132), .D1(n20_adj_4636), .CIN(n15692), .COUT(n15693), 
          .S0(d8_71__N_1603_adj_5707[52]), .S1(d8_71__N_1603_adj_5707[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_17 (.A0(d7_adj_5680[50]), .B0(cout_adj_5303), 
          .C0(n141), .D0(n23_adj_4633), .A1(d7_adj_5680[51]), .B1(cout_adj_5303), 
          .C1(n138), .D1(n22_adj_4634), .CIN(n15691), .COUT(n15692), 
          .S0(d8_71__N_1603_adj_5707[50]), .S1(d8_71__N_1603_adj_5707[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_15 (.A0(d7_adj_5680[48]), .B0(cout_adj_5303), 
          .C0(n147), .D0(n25_adj_4631), .A1(d7_adj_5680[49]), .B1(cout_adj_5303), 
          .C1(n144), .D1(n24_adj_4632), .CIN(n15690), .COUT(n15691), 
          .S0(d8_71__N_1603_adj_5707[48]), .S1(d8_71__N_1603_adj_5707[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_13 (.A0(d7_adj_5680[46]), .B0(cout_adj_5303), 
          .C0(n153), .D0(n27_adj_4629), .A1(d7_adj_5680[47]), .B1(cout_adj_5303), 
          .C1(n150), .D1(n26_adj_4630), .CIN(n15689), .COUT(n15690), 
          .S0(d8_71__N_1603_adj_5707[46]), .S1(d8_71__N_1603_adj_5707[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_11 (.A0(d7_adj_5680[44]), .B0(cout_adj_5303), 
          .C0(n159), .D0(n29_adj_4627), .A1(d7_adj_5680[45]), .B1(cout_adj_5303), 
          .C1(n156), .D1(n28_adj_4628), .CIN(n15688), .COUT(n15689), 
          .S0(d8_71__N_1603_adj_5707[44]), .S1(d8_71__N_1603_adj_5707[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_9 (.A0(d7_adj_5680[42]), .B0(cout_adj_5303), 
          .C0(n165), .D0(n31_adj_4624), .A1(d7_adj_5680[43]), .B1(cout_adj_5303), 
          .C1(n162), .D1(n30_adj_4626), .CIN(n15687), .COUT(n15688), 
          .S0(d8_71__N_1603_adj_5707[42]), .S1(d8_71__N_1603_adj_5707[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_7 (.A0(d7_adj_5680[40]), .B0(cout_adj_5303), 
          .C0(n171), .D0(n33_adj_4622), .A1(d7_adj_5680[41]), .B1(cout_adj_5303), 
          .C1(n168), .D1(n32_adj_4623), .CIN(n15686), .COUT(n15687), 
          .S0(d8_71__N_1603_adj_5707[40]), .S1(d8_71__N_1603_adj_5707[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_5 (.A0(d7_adj_5680[38]), .B0(cout_adj_5303), 
          .C0(n177), .D0(n35_adj_4620), .A1(d7_adj_5680[39]), .B1(cout_adj_5303), 
          .C1(n174), .D1(n34_adj_4621), .CIN(n15685), .COUT(n15686), 
          .S0(d8_71__N_1603_adj_5707[38]), .S1(d8_71__N_1603_adj_5707[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_3 (.A0(d7_adj_5680[36]), .B0(cout_adj_5303), 
          .C0(n183), .D0(n37_adj_4618), .A1(d7_adj_5680[37]), .B1(cout_adj_5303), 
          .C1(n180), .D1(n36_adj_4619), .CIN(n15684), .COUT(n15685), 
          .S0(d8_71__N_1603_adj_5707[36]), .S1(d8_71__N_1603_adj_5707[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5303), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15684));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1475_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1475_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15680), .S0(cout_adj_5088));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1424_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1424_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_36 (.A0(d5[34]), .B0(d4[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[35]), .B1(d4[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15679), .COUT(n15680), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_34 (.A0(d5[32]), .B0(d4[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[33]), .B1(d4[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15678), .COUT(n15679), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_32 (.A0(d5[30]), .B0(d4[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[31]), .B1(d4[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15677), .COUT(n15678), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_30 (.A0(d5[28]), .B0(d4[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[29]), .B1(d4[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15676), .COUT(n15677), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_28 (.A0(d5[26]), .B0(d4[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[27]), .B1(d4[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15675), .COUT(n15676), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_26 (.A0(d5[24]), .B0(d4[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[25]), .B1(d4[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15674), .COUT(n15675), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_24 (.A0(d5[22]), .B0(d4[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[23]), .B1(d4[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15673), .COUT(n15674), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_22 (.A0(d5[20]), .B0(d4[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[21]), .B1(d4[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15672), .COUT(n15673), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_20 (.A0(d5[18]), .B0(d4[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[19]), .B1(d4[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15671), .COUT(n15672), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_18 (.A0(d5[16]), .B0(d4[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[17]), .B1(d4[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15670), .COUT(n15671), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_16 (.A0(d5[14]), .B0(d4[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[15]), .B1(d4[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15669), .COUT(n15670), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_14 (.A0(d5[12]), .B0(d4[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[13]), .B1(d4[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15668), .COUT(n15669), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_12 (.A0(d5[10]), .B0(d4[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[11]), .B1(d4[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15667), .COUT(n15668), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_10 (.A0(d5[8]), .B0(d4[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[9]), .B1(d4[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15666), .COUT(n15667), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_8 (.A0(d5[6]), .B0(d4[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[7]), .B1(d4[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15665), 
          .COUT(n15666), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_6 (.A0(d5[4]), .B0(d4[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[5]), .B1(d4[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15664), 
          .COUT(n15665), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_4 (.A0(d5[2]), .B0(d4[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[3]), .B1(d4[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15663), 
          .COUT(n15664), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_2 (.A0(d5[0]), .B0(d4[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[1]), .B1(d4[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15663), 
          .S1(d5_71__N_706[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1424_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15661), .S0(cout_adj_5089));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1427_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1427_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_36 (.A0(d1_adj_5673[34]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[35]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15660), .COUT(n15661), .S0(d1_71__N_418_adj_5689[34]), 
          .S1(d1_71__N_418_adj_5689[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_34 (.A0(d1_adj_5673[32]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[33]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15659), .COUT(n15660), .S0(d1_71__N_418_adj_5689[32]), 
          .S1(d1_71__N_418_adj_5689[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_32 (.A0(d1_adj_5673[30]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[31]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15658), .COUT(n15659), .S0(d1_71__N_418_adj_5689[30]), 
          .S1(d1_71__N_418_adj_5689[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_30 (.A0(d1_adj_5673[28]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[29]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15657), .COUT(n15658), .S0(d1_71__N_418_adj_5689[28]), 
          .S1(d1_71__N_418_adj_5689[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_28 (.A0(d1_adj_5673[26]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[27]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15656), .COUT(n15657), .S0(d1_71__N_418_adj_5689[26]), 
          .S1(d1_71__N_418_adj_5689[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_26 (.A0(d1_adj_5673[24]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[25]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15655), .COUT(n15656), .S0(d1_71__N_418_adj_5689[24]), 
          .S1(d1_71__N_418_adj_5689[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_24 (.A0(d1_adj_5673[22]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[23]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15654), .COUT(n15655), .S0(d1_71__N_418_adj_5689[22]), 
          .S1(d1_71__N_418_adj_5689[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_22 (.A0(d1_adj_5673[20]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[21]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15653), .COUT(n15654), .S0(d1_71__N_418_adj_5689[20]), 
          .S1(d1_71__N_418_adj_5689[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_20 (.A0(d1_adj_5673[18]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[19]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15652), .COUT(n15653), .S0(d1_71__N_418_adj_5689[18]), 
          .S1(d1_71__N_418_adj_5689[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_18 (.A0(d1_adj_5673[16]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[17]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15651), .COUT(n15652), .S0(d1_71__N_418_adj_5689[16]), 
          .S1(d1_71__N_418_adj_5689[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_16 (.A0(d1_adj_5673[14]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[15]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15650), .COUT(n15651), .S0(d1_71__N_418_adj_5689[14]), 
          .S1(d1_71__N_418_adj_5689[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_14 (.A0(d1_adj_5673[12]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[13]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15649), .COUT(n15650), .S0(d1_71__N_418_adj_5689[12]), 
          .S1(d1_71__N_418_adj_5689[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_12 (.A0(d1_adj_5673[10]), .B0(MixerOutCos[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[11]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15648), .COUT(n15649), .S0(d1_71__N_418_adj_5689[10]), 
          .S1(d1_71__N_418_adj_5689[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_10 (.A0(d1_adj_5673[8]), .B0(MixerOutCos[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[9]), .B1(MixerOutCos[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15647), .COUT(n15648), .S0(d1_71__N_418_adj_5689[8]), 
          .S1(d1_71__N_418_adj_5689[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_8 (.A0(d1_adj_5673[6]), .B0(MixerOutCos[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[7]), .B1(MixerOutCos[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15646), .COUT(n15647), .S0(d1_71__N_418_adj_5689[6]), 
          .S1(d1_71__N_418_adj_5689[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_6 (.A0(d1_adj_5673[4]), .B0(MixerOutCos[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[5]), .B1(MixerOutCos[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15645), .COUT(n15646), .S0(d1_71__N_418_adj_5689[4]), 
          .S1(d1_71__N_418_adj_5689[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_4 (.A0(d1_adj_5673[2]), .B0(MixerOutCos[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[3]), .B1(MixerOutCos[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15644), .COUT(n15645), .S0(d1_71__N_418_adj_5689[2]), 
          .S1(d1_71__N_418_adj_5689[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_2 (.A0(d1_adj_5673[0]), .B0(MixerOutCos[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[1]), .B1(MixerOutCos[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15644), .S1(d1_71__N_418_adj_5689[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1427_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15642), .S0(n36_adj_5090));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1430_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15641), .COUT(n15642), .S0(n42), .S1(n39));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15640), .COUT(n15641), .S0(n48), .S1(n45));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15639), .COUT(n15640), .S0(n54), .S1(n51));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15638), .COUT(n15639), .S0(n60), .S1(n57));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15637), .COUT(n15638), .S0(n66_adj_5092), .S1(n63_adj_5091));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15636), .COUT(n15637), .S0(n72), .S1(n69));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15635), .COUT(n15636), .S0(n78_adj_5093), .S1(n75));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15635), .S1(n81_adj_5094));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1430_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1430_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_38 (.A0(d1[71]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15634), .S0(n78_adj_5095));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1553_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_36 (.A0(d1[69]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[70]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15633), .COUT(n15634), .S0(n84_adj_5097), 
          .S1(n81_adj_5096));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_34 (.A0(d1[67]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[68]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15632), .COUT(n15633), .S0(n90_adj_5099), 
          .S1(n87_adj_5098));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_32 (.A0(d1[65]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[66]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15631), .COUT(n15632), .S0(n96_adj_5101), 
          .S1(n93_adj_5100));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_30 (.A0(d1[63]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[64]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15630), .COUT(n15631), .S0(n102_adj_5103), 
          .S1(n99_adj_5102));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_28 (.A0(d1[61]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[62]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15629), .COUT(n15630), .S0(n108_adj_5105), 
          .S1(n105_adj_5104));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_26 (.A0(d1[59]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[60]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15628), .COUT(n15629), .S0(n114_adj_5107), 
          .S1(n111_adj_5106));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_24 (.A0(d1[57]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[58]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15627), .COUT(n15628), .S0(n120_adj_5109), 
          .S1(n117_adj_5108));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_22 (.A0(d1[55]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[56]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15626), .COUT(n15627), .S0(n126_adj_5111), 
          .S1(n123_adj_5110));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_20 (.A0(d1[53]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[54]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15625), .COUT(n15626), .S0(n132_adj_5113), 
          .S1(n129_adj_5112));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_18 (.A0(d1[51]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[52]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15624), .COUT(n15625), .S0(n138_adj_5115), 
          .S1(n135_adj_5114));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_16 (.A0(d1[49]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[50]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15623), .COUT(n15624), .S0(n144_adj_5117), 
          .S1(n141_adj_5116));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_14 (.A0(d1[47]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[48]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15622), .COUT(n15623), .S0(n150_adj_5119), 
          .S1(n147_adj_5118));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_12 (.A0(d1[45]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[46]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15621), .COUT(n15622), .S0(n156_adj_5121), 
          .S1(n153_adj_5120));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_10 (.A0(d1[43]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[44]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15620), .COUT(n15621), .S0(n162_adj_5123), 
          .S1(n159_adj_5122));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_8 (.A0(d1[41]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[42]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15619), .COUT(n15620), .S0(n168_adj_5125), 
          .S1(n165_adj_5124));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_6 (.A0(d1[39]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[40]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15618), .COUT(n15619), .S0(n174_adj_5127), 
          .S1(n171_adj_5126));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_4 (.A0(d1[37]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[38]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15617), .COUT(n15618), .S0(n180_adj_5129), 
          .S1(n177_adj_5128));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[36]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15617), .S1(n183_adj_5130));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1553_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1553_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15616), .S0(cout));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1415_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1415_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_36 (.A0(d2[34]), .B0(d1[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[35]), .B1(d1[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15615), .COUT(n15616), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_34 (.A0(d2[32]), .B0(d1[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[33]), .B1(d1[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15614), .COUT(n15615), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_32 (.A0(d2[30]), .B0(d1[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[31]), .B1(d1[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15613), .COUT(n15614), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_30 (.A0(d2[28]), .B0(d1[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[29]), .B1(d1[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15612), .COUT(n15613), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_30.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i3 (.D(n120_adj_5189), .CK(CIC1_out_clkSin), .Q(ISquare[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i3.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i4 (.D(n117_adj_5188), .CK(CIC1_out_clkSin), .Q(ISquare[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i4.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i5 (.D(n114_adj_5187), .CK(CIC1_out_clkSin), .Q(ISquare[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i5.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i6 (.D(n111_adj_5186), .CK(CIC1_out_clkSin), .Q(ISquare[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i6.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i7 (.D(n108_adj_5185), .CK(CIC1_out_clkSin), .Q(ISquare[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i7.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i8 (.D(n105_adj_5184), .CK(CIC1_out_clkSin), .Q(ISquare[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i8.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i9 (.D(n102_adj_5183), .CK(CIC1_out_clkSin), .Q(ISquare[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i9.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i10 (.D(n99_adj_5182), .CK(CIC1_out_clkSin), .Q(ISquare[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i10.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i11 (.D(n96_adj_5181), .CK(CIC1_out_clkSin), .Q(ISquare[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i11.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i12 (.D(n93_adj_5180), .CK(CIC1_out_clkSin), .Q(ISquare[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i12.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i13 (.D(n90_adj_5179), .CK(CIC1_out_clkSin), .Q(ISquare[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i13.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i14 (.D(n87_adj_5178), .CK(CIC1_out_clkSin), .Q(ISquare[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i14.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i15 (.D(n84_adj_5177), .CK(CIC1_out_clkSin), .Q(ISquare[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i15.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i16 (.D(n81_adj_5176), .CK(CIC1_out_clkSin), .Q(ISquare[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i16.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i17 (.D(n78_adj_5175), .CK(CIC1_out_clkSin), .Q(ISquare[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i17.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i18 (.D(n75_adj_5174), .CK(CIC1_out_clkSin), .Q(ISquare[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i18.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i19 (.D(n72_adj_5173), .CK(CIC1_out_clkSin), .Q(ISquare[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i19.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i20 (.D(n69_adj_5172), .CK(CIC1_out_clkSin), .Q(ISquare[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i20.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i21 (.D(n66_adj_5171), .CK(CIC1_out_clkSin), .Q(ISquare[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i21.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i22 (.D(n63_adj_5170), .CK(CIC1_out_clkSin), .Q(ISquare[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i22.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i23 (.D(n60_adj_5169), .CK(CIC1_out_clkSin), .Q(ISquare[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i23.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i24 (.D(n57_adj_5168), .CK(CIC1_out_clkSin), .Q(ISquare[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i24.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i25 (.D(n54_adj_5167), .CK(CIC1_out_clkSin), .Q(ISquare[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i25.GSR = "ENABLED";
    CCU2C _add_1_1415_add_4_28 (.A0(d2[26]), .B0(d1[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[27]), .B1(d1[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15611), .COUT(n15612), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_26 (.A0(d2[24]), .B0(d1[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[25]), .B1(d1[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15610), .COUT(n15611), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_24 (.A0(d2[22]), .B0(d1[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[23]), .B1(d1[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15609), .COUT(n15610), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_22 (.A0(d2[20]), .B0(d1[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[21]), .B1(d1[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15608), .COUT(n15609), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_20 (.A0(d2[18]), .B0(d1[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[19]), .B1(d1[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15607), .COUT(n15608), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_18 (.A0(d2[16]), .B0(d1[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[17]), .B1(d1[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15606), .COUT(n15607), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_16 (.A0(d2[14]), .B0(d1[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[15]), .B1(d1[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15605), .COUT(n15606), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_14 (.A0(d2[12]), .B0(d1[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[13]), .B1(d1[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15604), .COUT(n15605), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_12 (.A0(d2[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[11]), .B1(d1[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15603), .COUT(n15604), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_10 (.A0(d2[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[9]), .B1(d1[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15602), .COUT(n15603), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_8 (.A0(d2[6]), .B0(d1[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[7]), .B1(d1[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15601), 
          .COUT(n15602), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_6 (.A0(d2[4]), .B0(d1[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[5]), .B1(d1[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15600), 
          .COUT(n15601), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_4 (.A0(d2[2]), .B0(d1[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[3]), .B1(d1[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15599), 
          .COUT(n15600), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_2 (.A0(d2[0]), .B0(d1[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[1]), .B1(d1[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15599), 
          .S1(d2_71__N_490[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1415_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_38 (.A0(d_d8[35]), .B0(d8[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15597), .S0(d9_71__N_1675[35]), .S1(cout_adj_4998));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1652_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_36 (.A0(d_d8[33]), .B0(d8[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[34]), .B1(d8[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15596), .COUT(n15597), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_34 (.A0(d_d8[31]), .B0(d8[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[32]), .B1(d8[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15595), .COUT(n15596), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_32 (.A0(d_d8[29]), .B0(d8[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[30]), .B1(d8[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15594), .COUT(n15595), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_30 (.A0(d_d8[27]), .B0(d8[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[28]), .B1(d8[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15593), .COUT(n15594), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_28 (.A0(d_d8[25]), .B0(d8[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[26]), .B1(d8[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15592), .COUT(n15593), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_26 (.A0(d_d8[23]), .B0(d8[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[24]), .B1(d8[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15591), .COUT(n15592), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_24 (.A0(d_d8[21]), .B0(d8[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[22]), .B1(d8[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15590), .COUT(n15591), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_22 (.A0(d_d8[19]), .B0(d8[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[20]), .B1(d8[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15589), .COUT(n15590), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_20 (.A0(d_d8[17]), .B0(d8[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[18]), .B1(d8[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15588), .COUT(n15589), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_18 (.A0(d_d8[15]), .B0(d8[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[16]), .B1(d8[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15587), .COUT(n15588), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_16 (.A0(d_d8[13]), .B0(d8[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[14]), .B1(d8[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15586), .COUT(n15587), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_14 (.A0(d_d8[11]), .B0(d8[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[12]), .B1(d8[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15585), .COUT(n15586), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_12 (.A0(d_d8[9]), .B0(d8[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[10]), .B1(d8[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15584), .COUT(n15585), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_10 (.A0(d_d8[7]), .B0(d8[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[8]), .B1(d8[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15583), .COUT(n15584), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_8 (.A0(d_d8[5]), .B0(d8[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[6]), .B1(d8[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15582), .COUT(n15583), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_6 (.A0(d_d8[3]), .B0(d8[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[4]), .B1(d8[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15581), .COUT(n15582), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_4 (.A0(d_d8[1]), .B0(d8[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[2]), .B1(d8[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15580), .COUT(n15581), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1652_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[0]), .B1(d8[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15580), .S1(d9_71__N_1675[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1652_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1652_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1652_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15579), .S0(cout_adj_4736));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1418_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1418_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_36 (.A0(d3[34]), .B0(d2[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[35]), .B1(d2[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15578), .COUT(n15579), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_34 (.A0(d3[32]), .B0(d2[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[33]), .B1(d2[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15577), .COUT(n15578), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_32 (.A0(d3[30]), .B0(d2[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[31]), .B1(d2[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15576), .COUT(n15577), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_30 (.A0(d3[28]), .B0(d2[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[29]), .B1(d2[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15575), .COUT(n15576), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_28 (.A0(d3[26]), .B0(d2[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[27]), .B1(d2[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15574), .COUT(n15575), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_26 (.A0(d3[24]), .B0(d2[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[25]), .B1(d2[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15573), .COUT(n15574), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_24 (.A0(d3[22]), .B0(d2[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[23]), .B1(d2[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15572), .COUT(n15573), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_22 (.A0(d3[20]), .B0(d2[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[21]), .B1(d2[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15571), .COUT(n15572), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_20 (.A0(d3[18]), .B0(d2[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[19]), .B1(d2[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15570), .COUT(n15571), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_18 (.A0(d3[16]), .B0(d2[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[17]), .B1(d2[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15569), .COUT(n15570), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_16 (.A0(d3[14]), .B0(d2[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[15]), .B1(d2[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15568), .COUT(n15569), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_14 (.A0(d3[12]), .B0(d2[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[13]), .B1(d2[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15567), .COUT(n15568), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_12 (.A0(d3[10]), .B0(d2[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[11]), .B1(d2[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15566), .COUT(n15567), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_10 (.A0(d3[8]), .B0(d2[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[9]), .B1(d2[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15565), .COUT(n15566), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_8 (.A0(d3[6]), .B0(d2[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[7]), .B1(d2[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15564), 
          .COUT(n15565), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_6 (.A0(d3[4]), .B0(d2[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[5]), .B1(d2[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15563), 
          .COUT(n15564), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_4 (.A0(d3[2]), .B0(d2[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[3]), .B1(d2[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15562), 
          .COUT(n15563), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_2 (.A0(d3[0]), .B0(d2[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[1]), .B1(d2[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15562), 
          .S1(d3_71__N_562[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1418_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_2.INJECT1_1 = "NO";
    LUT4 i3172_2_lut (.A(led_c_4), .B(n2845), .Z(n3715)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3172_2_lut.init = 16'h4444;
    CCU2C _add_1_1580_add_4_38 (.A0(d5_adj_5677[71]), .B0(d4_adj_5676[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15560), .S0(n78_adj_4837));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1580_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_36 (.A0(d5_adj_5677[69]), .B0(d4_adj_5676[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[70]), .B1(d4_adj_5676[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15559), .COUT(n15560), .S0(n84_adj_4839), 
          .S1(n81_adj_4838));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_34 (.A0(d5_adj_5677[67]), .B0(d4_adj_5676[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[68]), .B1(d4_adj_5676[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15558), .COUT(n15559), .S0(n90_adj_4841), 
          .S1(n87_adj_4840));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_32 (.A0(d5_adj_5677[65]), .B0(d4_adj_5676[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[66]), .B1(d4_adj_5676[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15557), .COUT(n15558), .S0(n96_adj_4843), 
          .S1(n93_adj_4842));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_30 (.A0(d5_adj_5677[63]), .B0(d4_adj_5676[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[64]), .B1(d4_adj_5676[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15556), .COUT(n15557), .S0(n102_adj_4845), 
          .S1(n99_adj_4844));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_28 (.A0(d5_adj_5677[61]), .B0(d4_adj_5676[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[62]), .B1(d4_adj_5676[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15555), .COUT(n15556), .S0(n108_adj_4847), 
          .S1(n105_adj_4846));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_26 (.A0(d5_adj_5677[59]), .B0(d4_adj_5676[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[60]), .B1(d4_adj_5676[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15554), .COUT(n15555), .S0(n114_adj_4849), 
          .S1(n111_adj_4848));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_24 (.A0(d5_adj_5677[57]), .B0(d4_adj_5676[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[58]), .B1(d4_adj_5676[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15553), .COUT(n15554), .S0(n120_adj_4851), 
          .S1(n117_adj_4850));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_22 (.A0(d5_adj_5677[55]), .B0(d4_adj_5676[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[56]), .B1(d4_adj_5676[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15552), .COUT(n15553), .S0(n126_adj_4853), 
          .S1(n123_adj_4852));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_20 (.A0(d5_adj_5677[53]), .B0(d4_adj_5676[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[54]), .B1(d4_adj_5676[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15551), .COUT(n15552), .S0(n132_adj_4855), 
          .S1(n129_adj_4854));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_18 (.A0(d5_adj_5677[51]), .B0(d4_adj_5676[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[52]), .B1(d4_adj_5676[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15550), .COUT(n15551), .S0(n138_adj_4857), 
          .S1(n135_adj_4856));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_16 (.A0(d5_adj_5677[49]), .B0(d4_adj_5676[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[50]), .B1(d4_adj_5676[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15549), .COUT(n15550), .S0(n144_adj_4859), 
          .S1(n141_adj_4858));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_14 (.A0(d5_adj_5677[47]), .B0(d4_adj_5676[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[48]), .B1(d4_adj_5676[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15548), .COUT(n15549), .S0(n150_adj_4861), 
          .S1(n147_adj_4860));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_12 (.A0(d5_adj_5677[45]), .B0(d4_adj_5676[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[46]), .B1(d4_adj_5676[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15547), .COUT(n15548), .S0(n156_adj_4863), 
          .S1(n153_adj_4862));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_10 (.A0(d5_adj_5677[43]), .B0(d4_adj_5676[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[44]), .B1(d4_adj_5676[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15546), .COUT(n15547), .S0(n162_adj_4865), 
          .S1(n159_adj_4864));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_8 (.A0(d5_adj_5677[41]), .B0(d4_adj_5676[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[42]), .B1(d4_adj_5676[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15545), .COUT(n15546), .S0(n168_adj_4867), 
          .S1(n165_adj_4866));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_6 (.A0(d5_adj_5677[39]), .B0(d4_adj_5676[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[40]), .B1(d4_adj_5676[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15544), .COUT(n15545), .S0(n174_adj_4869), 
          .S1(n171_adj_4868));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_4 (.A0(d5_adj_5677[37]), .B0(d4_adj_5676[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5677[38]), .B1(d4_adj_5676[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15543), .COUT(n15544), .S0(n180_adj_4871), 
          .S1(n177_adj_4870));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1580_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5_adj_5677[36]), .B1(d4_adj_5676[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15543), .S1(n183_adj_4872));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1580_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1580_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1580_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_37 (.A0(d8_adj_5682[70]), .B0(cout_adj_5230), 
          .C0(n81_adj_4874), .D0(n3_adj_4615), .A1(d8_adj_5682[71]), .B1(cout_adj_5230), 
          .C1(n78_adj_4873), .D1(n2_adj_4616), .CIN(n15541), .S0(d9_71__N_1675_adj_5708[70]), 
          .S1(d9_71__N_1675_adj_5708[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_35 (.A0(d8_adj_5682[68]), .B0(cout_adj_5230), 
          .C0(n87_adj_4876), .D0(n5_adj_4613), .A1(d8_adj_5682[69]), .B1(cout_adj_5230), 
          .C1(n84_adj_4875), .D1(n4_adj_4614), .CIN(n15540), .COUT(n15541), 
          .S0(d9_71__N_1675_adj_5708[68]), .S1(d9_71__N_1675_adj_5708[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_33 (.A0(d8_adj_5682[66]), .B0(cout_adj_5230), 
          .C0(n93_adj_4878), .D0(n7_adj_4611), .A1(d8_adj_5682[67]), .B1(cout_adj_5230), 
          .C1(n90_adj_4877), .D1(n6_adj_4612), .CIN(n15539), .COUT(n15540), 
          .S0(d9_71__N_1675_adj_5708[66]), .S1(d9_71__N_1675_adj_5708[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_31 (.A0(d8_adj_5682[64]), .B0(cout_adj_5230), 
          .C0(n99_adj_4880), .D0(n9_adj_4609), .A1(d8_adj_5682[65]), .B1(cout_adj_5230), 
          .C1(n96_adj_4879), .D1(n8_adj_4610), .CIN(n15538), .COUT(n15539), 
          .S0(d9_71__N_1675_adj_5708[64]), .S1(d9_71__N_1675_adj_5708[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_29 (.A0(d8_adj_5682[62]), .B0(cout_adj_5230), 
          .C0(n105_adj_4882), .D0(n11_adj_4607), .A1(d8_adj_5682[63]), 
          .B1(cout_adj_5230), .C1(n102_adj_4881), .D1(n10_adj_4608), .CIN(n15537), 
          .COUT(n15538), .S0(d9_71__N_1675_adj_5708[62]), .S1(d9_71__N_1675_adj_5708[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_27 (.A0(d8_adj_5682[60]), .B0(cout_adj_5230), 
          .C0(n111_adj_4884), .D0(n13_adj_4605), .A1(d8_adj_5682[61]), 
          .B1(cout_adj_5230), .C1(n108_adj_4883), .D1(n12_adj_4606), .CIN(n15536), 
          .COUT(n15537), .S0(d9_71__N_1675_adj_5708[60]), .S1(d9_71__N_1675_adj_5708[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_25 (.A0(d8_adj_5682[58]), .B0(cout_adj_5230), 
          .C0(n117_adj_4886), .D0(n15_adj_4603), .A1(d8_adj_5682[59]), 
          .B1(cout_adj_5230), .C1(n114_adj_4885), .D1(n14_adj_4604), .CIN(n15535), 
          .COUT(n15536), .S0(d9_71__N_1675_adj_5708[58]), .S1(d9_71__N_1675_adj_5708[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_23 (.A0(d8_adj_5682[56]), .B0(cout_adj_5230), 
          .C0(n123_adj_4888), .D0(n17_adj_4601), .A1(d8_adj_5682[57]), 
          .B1(cout_adj_5230), .C1(n120_adj_4887), .D1(n16_adj_4602), .CIN(n15534), 
          .COUT(n15535), .S0(d9_71__N_1675_adj_5708[56]), .S1(d9_71__N_1675_adj_5708[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_21 (.A0(d8_adj_5682[54]), .B0(cout_adj_5230), 
          .C0(n129_adj_4890), .D0(n19_adj_4599), .A1(d8_adj_5682[55]), 
          .B1(cout_adj_5230), .C1(n126_adj_4889), .D1(n18_adj_4600), .CIN(n15533), 
          .COUT(n15534), .S0(d9_71__N_1675_adj_5708[54]), .S1(d9_71__N_1675_adj_5708[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_19 (.A0(d8_adj_5682[52]), .B0(cout_adj_5230), 
          .C0(n135_adj_4892), .D0(n21_adj_4597), .A1(d8_adj_5682[53]), 
          .B1(cout_adj_5230), .C1(n132_adj_4891), .D1(n20_adj_4598), .CIN(n15532), 
          .COUT(n15533), .S0(d9_71__N_1675_adj_5708[52]), .S1(d9_71__N_1675_adj_5708[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_17 (.A0(d8_adj_5682[50]), .B0(cout_adj_5230), 
          .C0(n141_adj_4894), .D0(n23_adj_4595), .A1(d8_adj_5682[51]), 
          .B1(cout_adj_5230), .C1(n138_adj_4893), .D1(n22_adj_4596), .CIN(n15531), 
          .COUT(n15532), .S0(d9_71__N_1675_adj_5708[50]), .S1(d9_71__N_1675_adj_5708[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_15 (.A0(d8_adj_5682[48]), .B0(cout_adj_5230), 
          .C0(n147_adj_4896), .D0(n25_adj_4593), .A1(d8_adj_5682[49]), 
          .B1(cout_adj_5230), .C1(n144_adj_4895), .D1(n24_adj_4594), .CIN(n15530), 
          .COUT(n15531), .S0(d9_71__N_1675_adj_5708[48]), .S1(d9_71__N_1675_adj_5708[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_13 (.A0(d8_adj_5682[46]), .B0(cout_adj_5230), 
          .C0(n153_adj_4898), .D0(n27_adj_4588), .A1(d8_adj_5682[47]), 
          .B1(cout_adj_5230), .C1(n150_adj_4897), .D1(n26_adj_4589), .CIN(n15529), 
          .COUT(n15530), .S0(d9_71__N_1675_adj_5708[46]), .S1(d9_71__N_1675_adj_5708[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_11 (.A0(d8_adj_5682[44]), .B0(cout_adj_5230), 
          .C0(n159_adj_4900), .D0(n29_adj_4586), .A1(d8_adj_5682[45]), 
          .B1(cout_adj_5230), .C1(n156_adj_4899), .D1(n28_adj_4587), .CIN(n15528), 
          .COUT(n15529), .S0(d9_71__N_1675_adj_5708[44]), .S1(d9_71__N_1675_adj_5708[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_9 (.A0(d8_adj_5682[42]), .B0(cout_adj_5230), 
          .C0(n165_adj_4902), .D0(n31_adj_4584), .A1(d8_adj_5682[43]), 
          .B1(cout_adj_5230), .C1(n162_adj_4901), .D1(n30_adj_4585), .CIN(n15527), 
          .COUT(n15528), .S0(d9_71__N_1675_adj_5708[42]), .S1(d9_71__N_1675_adj_5708[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_7 (.A0(d8_adj_5682[40]), .B0(cout_adj_5230), 
          .C0(n171_adj_4904), .D0(n33_adj_4582), .A1(d8_adj_5682[41]), 
          .B1(cout_adj_5230), .C1(n168_adj_4903), .D1(n32_adj_4583), .CIN(n15526), 
          .COUT(n15527), .S0(d9_71__N_1675_adj_5708[40]), .S1(d9_71__N_1675_adj_5708[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_5 (.A0(d8_adj_5682[38]), .B0(cout_adj_5230), 
          .C0(n177_adj_4906), .D0(n35_adj_4580), .A1(d8_adj_5682[39]), 
          .B1(cout_adj_5230), .C1(n174_adj_4905), .D1(n34_adj_4581), .CIN(n15525), 
          .COUT(n15526), .S0(d9_71__N_1675_adj_5708[38]), .S1(d9_71__N_1675_adj_5708[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_3 (.A0(d8_adj_5682[36]), .B0(cout_adj_5230), 
          .C0(n183_adj_4908), .D0(n37_adj_4578), .A1(d8_adj_5682[37]), 
          .B1(cout_adj_5230), .C1(n180_adj_4907), .D1(n36_adj_4579), .CIN(n15524), 
          .COUT(n15525), .S0(d9_71__N_1675_adj_5708[36]), .S1(d9_71__N_1675_adj_5708[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5230), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15524));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1472_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1472_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15520), .S0(cout_adj_5663));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1406_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1406_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_36 (.A0(d1[34]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[35]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15519), .COUT(n15520), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_34 (.A0(d1[32]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[33]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15518), .COUT(n15519), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_32 (.A0(d1[30]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[31]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15517), .COUT(n15518), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_30 (.A0(d1[28]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[29]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15516), .COUT(n15517), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_28 (.A0(d1[26]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[27]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15515), .COUT(n15516), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_26 (.A0(d1[24]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[25]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15514), .COUT(n15515), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_24 (.A0(d1[22]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[23]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15513), .COUT(n15514), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_22 (.A0(d1[20]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[21]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15512), .COUT(n15513), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_20 (.A0(d1[18]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[19]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15511), .COUT(n15512), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_18 (.A0(d1[16]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[17]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15510), .COUT(n15511), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_16 (.A0(d1[14]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[15]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15509), .COUT(n15510), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_14 (.A0(d1[12]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[13]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15508), .COUT(n15509), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_12 (.A0(d1[10]), .B0(MixerOutSin[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[11]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15507), .COUT(n15508), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_10 (.A0(d1[8]), .B0(MixerOutSin[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[9]), .B1(MixerOutSin[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15506), .COUT(n15507), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_8 (.A0(d1[6]), .B0(MixerOutSin[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[7]), .B1(MixerOutSin[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15505), .COUT(n15506), .S0(d1_71__N_418[6]), 
          .S1(d1_71__N_418[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_6 (.A0(d1[4]), .B0(MixerOutSin[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[5]), .B1(MixerOutSin[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15504), .COUT(n15505), .S0(d1_71__N_418[4]), 
          .S1(d1_71__N_418[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_4 (.A0(d1[2]), .B0(MixerOutSin[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[3]), .B1(MixerOutSin[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15503), .COUT(n15504), .S0(d1_71__N_418[2]), 
          .S1(d1_71__N_418[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_2 (.A0(d1[0]), .B0(MixerOutSin[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[1]), .B1(MixerOutSin[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15503), .S1(d1_71__N_418[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1406_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1406_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_38 (.A0(d3_adj_5675[71]), .B0(d2_adj_5674[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15501), .S0(n78_adj_5623));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1574_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_36 (.A0(d3_adj_5675[69]), .B0(d2_adj_5674[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[70]), .B1(d2_adj_5674[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15500), .COUT(n15501), .S0(n84_adj_5625), 
          .S1(n81_adj_5624));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_34 (.A0(d3_adj_5675[67]), .B0(d2_adj_5674[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[68]), .B1(d2_adj_5674[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15499), .COUT(n15500), .S0(n90_adj_5627), 
          .S1(n87_adj_5626));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_32 (.A0(d3_adj_5675[65]), .B0(d2_adj_5674[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[66]), .B1(d2_adj_5674[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15498), .COUT(n15499), .S0(n96_adj_5629), 
          .S1(n93_adj_5628));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_30 (.A0(d3_adj_5675[63]), .B0(d2_adj_5674[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[64]), .B1(d2_adj_5674[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15497), .COUT(n15498), .S0(n102_adj_5631), 
          .S1(n99_adj_5630));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_28 (.A0(d3_adj_5675[61]), .B0(d2_adj_5674[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[62]), .B1(d2_adj_5674[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15496), .COUT(n15497), .S0(n108_adj_5633), 
          .S1(n105_adj_5632));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_26 (.A0(d3_adj_5675[59]), .B0(d2_adj_5674[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[60]), .B1(d2_adj_5674[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15495), .COUT(n15496), .S0(n114_adj_5635), 
          .S1(n111_adj_5634));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_24 (.A0(d3_adj_5675[57]), .B0(d2_adj_5674[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[58]), .B1(d2_adj_5674[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15494), .COUT(n15495), .S0(n120_adj_5637), 
          .S1(n117_adj_5636));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_22 (.A0(d3_adj_5675[55]), .B0(d2_adj_5674[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[56]), .B1(d2_adj_5674[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15493), .COUT(n15494), .S0(n126_adj_5639), 
          .S1(n123_adj_5638));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_20 (.A0(d3_adj_5675[53]), .B0(d2_adj_5674[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[54]), .B1(d2_adj_5674[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15492), .COUT(n15493), .S0(n132_adj_5641), 
          .S1(n129_adj_5640));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_18 (.A0(d3_adj_5675[51]), .B0(d2_adj_5674[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[52]), .B1(d2_adj_5674[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15491), .COUT(n15492), .S0(n138_adj_5643), 
          .S1(n135_adj_5642));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_16 (.A0(d3_adj_5675[49]), .B0(d2_adj_5674[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[50]), .B1(d2_adj_5674[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15490), .COUT(n15491), .S0(n144_adj_5645), 
          .S1(n141_adj_5644));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_14 (.A0(d3_adj_5675[47]), .B0(d2_adj_5674[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[48]), .B1(d2_adj_5674[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15489), .COUT(n15490), .S0(n150_adj_5647), 
          .S1(n147_adj_5646));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_12 (.A0(d3_adj_5675[45]), .B0(d2_adj_5674[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[46]), .B1(d2_adj_5674[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15488), .COUT(n15489), .S0(n156_adj_5649), 
          .S1(n153_adj_5648));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_10 (.A0(d3_adj_5675[43]), .B0(d2_adj_5674[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[44]), .B1(d2_adj_5674[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15487), .COUT(n15488), .S0(n162_adj_5651), 
          .S1(n159_adj_5650));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_8 (.A0(d3_adj_5675[41]), .B0(d2_adj_5674[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[42]), .B1(d2_adj_5674[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15486), .COUT(n15487), .S0(n168_adj_5653), 
          .S1(n165_adj_5652));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_6 (.A0(d3_adj_5675[39]), .B0(d2_adj_5674[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[40]), .B1(d2_adj_5674[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15485), .COUT(n15486), .S0(n174_adj_5655), 
          .S1(n171_adj_5654));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_4 (.A0(d3_adj_5675[37]), .B0(d2_adj_5674[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5675[38]), .B1(d2_adj_5674[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15484), .COUT(n15485), .S0(n180_adj_5657), 
          .S1(n177_adj_5656));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3_adj_5675[36]), .B1(d2_adj_5674[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15484), .S1(n183_adj_5658));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(66[13:20])
    defparam _add_1_1574_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1574_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_37 (.A0(d_d9_adj_5685[71]), .B0(d9_adj_5684[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15483), .S0(n76_adj_5545));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1469_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_35 (.A0(d_d9_adj_5685[69]), .B0(d9_adj_5684[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[70]), .B1(d9_adj_5684[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15482), .COUT(n15483), .S0(n82_adj_5547), 
          .S1(n79_adj_5546));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_33 (.A0(d_d9_adj_5685[67]), .B0(d9_adj_5684[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[68]), .B1(d9_adj_5684[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15481), .COUT(n15482), .S0(n88_adj_5549), 
          .S1(n85_adj_5548));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_31 (.A0(d_d9_adj_5685[65]), .B0(d9_adj_5684[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[66]), .B1(d9_adj_5684[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15480), .COUT(n15481), .S0(n94_adj_5551), 
          .S1(n91_adj_5550));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_29 (.A0(d_d9_adj_5685[63]), .B0(d9_adj_5684[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[64]), .B1(d9_adj_5684[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15479), .COUT(n15480), .S0(n100_adj_5553), 
          .S1(n97_adj_5552));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_27 (.A0(d_d9_adj_5685[61]), .B0(d9_adj_5684[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[62]), .B1(d9_adj_5684[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15478), .COUT(n15479), .S0(n106_adj_5555), 
          .S1(n103_adj_5554));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_25 (.A0(d_d9_adj_5685[59]), .B0(d9_adj_5684[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[60]), .B1(d9_adj_5684[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15477), .COUT(n15478), .S0(n112_adj_5557), 
          .S1(n109_adj_5556));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_23 (.A0(d_d9_adj_5685[57]), .B0(d9_adj_5684[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[58]), .B1(d9_adj_5684[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15476), .COUT(n15477), .S0(n118_adj_5559), 
          .S1(n115_adj_5558));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_21 (.A0(d_d9_adj_5685[55]), .B0(d9_adj_5684[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[56]), .B1(d9_adj_5684[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15475), .COUT(n15476));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_19 (.A0(d_d9_adj_5685[53]), .B0(d9_adj_5684[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[54]), .B1(d9_adj_5684[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15474), .COUT(n15475));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_17 (.A0(d_d9_adj_5685[51]), .B0(d9_adj_5684[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[52]), .B1(d9_adj_5684[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15473), .COUT(n15474));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_15 (.A0(d_d9_adj_5685[49]), .B0(d9_adj_5684[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[50]), .B1(d9_adj_5684[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15472), .COUT(n15473));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_13 (.A0(d_d9_adj_5685[47]), .B0(d9_adj_5684[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[48]), .B1(d9_adj_5684[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15471), .COUT(n15472));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_11 (.A0(d_d9_adj_5685[45]), .B0(d9_adj_5684[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[46]), .B1(d9_adj_5684[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15470), .COUT(n15471));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_9 (.A0(d_d9_adj_5685[43]), .B0(d9_adj_5684[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[44]), .B1(d9_adj_5684[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15469), .COUT(n15470));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_7 (.A0(d_d9_adj_5685[41]), .B0(d9_adj_5684[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[42]), .B1(d9_adj_5684[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15468), .COUT(n15469));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_5 (.A0(d_d9_adj_5685[39]), .B0(d9_adj_5684[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[40]), .B1(d9_adj_5684[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15467), .COUT(n15468));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_3 (.A0(d_d9_adj_5685[37]), .B0(d9_adj_5684[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[38]), .B1(d9_adj_5684[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15466), .COUT(n15467));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5685[36]), .B1(d9_adj_5684[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15466));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1469_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_38 (.A0(d_d8_adj_5683[71]), .B0(d8_adj_5682[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15465), .S0(n78_adj_4873));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1634_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_36 (.A0(d_d8_adj_5683[69]), .B0(d8_adj_5682[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[70]), .B1(d8_adj_5682[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15464), .COUT(n15465), .S0(n84_adj_4875), 
          .S1(n81_adj_4874));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_34 (.A0(d_d8_adj_5683[67]), .B0(d8_adj_5682[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[68]), .B1(d8_adj_5682[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15463), .COUT(n15464), .S0(n90_adj_4877), 
          .S1(n87_adj_4876));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_32 (.A0(d_d8_adj_5683[65]), .B0(d8_adj_5682[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[66]), .B1(d8_adj_5682[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15462), .COUT(n15463), .S0(n96_adj_4879), 
          .S1(n93_adj_4878));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_30 (.A0(d_d8_adj_5683[63]), .B0(d8_adj_5682[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[64]), .B1(d8_adj_5682[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15461), .COUT(n15462), .S0(n102_adj_4881), 
          .S1(n99_adj_4880));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_28 (.A0(d_d8_adj_5683[61]), .B0(d8_adj_5682[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[62]), .B1(d8_adj_5682[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15460), .COUT(n15461), .S0(n108_adj_4883), 
          .S1(n105_adj_4882));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_26 (.A0(d_d8_adj_5683[59]), .B0(d8_adj_5682[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[60]), .B1(d8_adj_5682[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15459), .COUT(n15460), .S0(n114_adj_4885), 
          .S1(n111_adj_4884));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_24 (.A0(d_d8_adj_5683[57]), .B0(d8_adj_5682[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[58]), .B1(d8_adj_5682[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15458), .COUT(n15459), .S0(n120_adj_4887), 
          .S1(n117_adj_4886));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_22 (.A0(d_d8_adj_5683[55]), .B0(d8_adj_5682[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[56]), .B1(d8_adj_5682[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15457), .COUT(n15458), .S0(n126_adj_4889), 
          .S1(n123_adj_4888));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_20 (.A0(d_d8_adj_5683[53]), .B0(d8_adj_5682[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[54]), .B1(d8_adj_5682[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15456), .COUT(n15457), .S0(n132_adj_4891), 
          .S1(n129_adj_4890));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_18 (.A0(d_d8_adj_5683[51]), .B0(d8_adj_5682[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[52]), .B1(d8_adj_5682[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15455), .COUT(n15456), .S0(n138_adj_4893), 
          .S1(n135_adj_4892));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_16 (.A0(d_d8_adj_5683[49]), .B0(d8_adj_5682[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[50]), .B1(d8_adj_5682[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15454), .COUT(n15455), .S0(n144_adj_4895), 
          .S1(n141_adj_4894));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_14 (.A0(d_d8_adj_5683[47]), .B0(d8_adj_5682[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[48]), .B1(d8_adj_5682[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15453), .COUT(n15454), .S0(n150_adj_4897), 
          .S1(n147_adj_4896));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_12 (.A0(d_d8_adj_5683[45]), .B0(d8_adj_5682[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[46]), .B1(d8_adj_5682[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15452), .COUT(n15453), .S0(n156_adj_4899), 
          .S1(n153_adj_4898));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_10 (.A0(d_d8_adj_5683[43]), .B0(d8_adj_5682[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[44]), .B1(d8_adj_5682[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15451), .COUT(n15452), .S0(n162_adj_4901), 
          .S1(n159_adj_4900));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_8 (.A0(d_d8_adj_5683[41]), .B0(d8_adj_5682[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[42]), .B1(d8_adj_5682[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15450), .COUT(n15451), .S0(n168_adj_4903), 
          .S1(n165_adj_4902));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_6 (.A0(d_d8_adj_5683[39]), .B0(d8_adj_5682[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[40]), .B1(d8_adj_5682[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15449), .COUT(n15450), .S0(n174_adj_4905), 
          .S1(n171_adj_4904));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_4 (.A0(d_d8_adj_5683[37]), .B0(d8_adj_5682[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5683[38]), .B1(d8_adj_5682[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15448), .COUT(n15449), .S0(n180_adj_4907), 
          .S1(n177_adj_4906));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5683[36]), .B1(d8_adj_5682[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15448), .S1(n183_adj_4908));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1634_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1634_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_38 (.A0(d_d8[71]), .B0(d8[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15447), .S0(n78_adj_4999));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1583_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_36 (.A0(d_d8[69]), .B0(d8[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[70]), .B1(d8[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15446), .COUT(n15447), .S0(n84_adj_5001), .S1(n81_adj_5000));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_34 (.A0(d_d8[67]), .B0(d8[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[68]), .B1(d8[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15445), .COUT(n15446), .S0(n90_adj_5003), .S1(n87_adj_5002));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_32 (.A0(d_d8[65]), .B0(d8[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[66]), .B1(d8[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15444), .COUT(n15445), .S0(n96_adj_5005), .S1(n93_adj_5004));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_30 (.A0(d_d8[63]), .B0(d8[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[64]), .B1(d8[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15443), .COUT(n15444), .S0(n102_adj_5007), .S1(n99_adj_5006));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_28 (.A0(d_d8[61]), .B0(d8[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[62]), .B1(d8[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15442), .COUT(n15443), .S0(n108_adj_5009), .S1(n105_adj_5008));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_26 (.A0(d_d8[59]), .B0(d8[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[60]), .B1(d8[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15441), .COUT(n15442), .S0(n114_adj_5011), .S1(n111_adj_5010));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_24 (.A0(d_d8[57]), .B0(d8[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[58]), .B1(d8[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15440), .COUT(n15441), .S0(n120_adj_5013), .S1(n117_adj_5012));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_22 (.A0(d_d8[55]), .B0(d8[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[56]), .B1(d8[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15439), .COUT(n15440), .S0(n126_adj_5015), .S1(n123_adj_5014));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_20 (.A0(d_d8[53]), .B0(d8[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[54]), .B1(d8[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15438), .COUT(n15439), .S0(n132_adj_5017), .S1(n129_adj_5016));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_18 (.A0(d_d8[51]), .B0(d8[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[52]), .B1(d8[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15437), .COUT(n15438), .S0(n138_adj_5019), .S1(n135_adj_5018));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_16 (.A0(d_d8[49]), .B0(d8[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[50]), .B1(d8[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15436), .COUT(n15437), .S0(n144_adj_5021), .S1(n141_adj_5020));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_14 (.A0(d_d8[47]), .B0(d8[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[48]), .B1(d8[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15435), .COUT(n15436), .S0(n150_adj_5023), .S1(n147_adj_5022));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_12 (.A0(d_d8[45]), .B0(d8[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[46]), .B1(d8[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15434), .COUT(n15435), .S0(n156_adj_5025), .S1(n153_adj_5024));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_10 (.A0(d_d8[43]), .B0(d8[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[44]), .B1(d8[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15433), .COUT(n15434), .S0(n162_adj_5027), .S1(n159_adj_5026));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_8 (.A0(d_d8[41]), .B0(d8[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[42]), .B1(d8[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15432), .COUT(n15433), .S0(n168_adj_5029), .S1(n165_adj_5028));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_6 (.A0(d_d8[39]), .B0(d8[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[40]), .B1(d8[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15431), .COUT(n15432), .S0(n174_adj_5031), .S1(n171_adj_5030));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_4 (.A0(d_d8[37]), .B0(d8[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[38]), .B1(d8[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15430), .COUT(n15431), .S0(n180_adj_5033), .S1(n177_adj_5032));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[36]), .B1(d8[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15430), .S1(n183_adj_5034));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam _add_1_1583_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1583_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15429), .S0(cout_adj_5131));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1433_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1433_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_36 (.A0(d2_adj_5674[34]), .B0(d1_adj_5673[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[35]), .B1(d1_adj_5673[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15428), .COUT(n15429), .S0(d2_71__N_490_adj_5690[34]), 
          .S1(d2_71__N_490_adj_5690[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_34 (.A0(d2_adj_5674[32]), .B0(d1_adj_5673[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[33]), .B1(d1_adj_5673[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15427), .COUT(n15428), .S0(d2_71__N_490_adj_5690[32]), 
          .S1(d2_71__N_490_adj_5690[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_32 (.A0(d2_adj_5674[30]), .B0(d1_adj_5673[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[31]), .B1(d1_adj_5673[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15426), .COUT(n15427), .S0(d2_71__N_490_adj_5690[30]), 
          .S1(d2_71__N_490_adj_5690[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_30 (.A0(d2_adj_5674[28]), .B0(d1_adj_5673[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[29]), .B1(d1_adj_5673[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15425), .COUT(n15426), .S0(d2_71__N_490_adj_5690[28]), 
          .S1(d2_71__N_490_adj_5690[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_28 (.A0(d2_adj_5674[26]), .B0(d1_adj_5673[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[27]), .B1(d1_adj_5673[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15424), .COUT(n15425), .S0(d2_71__N_490_adj_5690[26]), 
          .S1(d2_71__N_490_adj_5690[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_26 (.A0(d2_adj_5674[24]), .B0(d1_adj_5673[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[25]), .B1(d1_adj_5673[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15423), .COUT(n15424), .S0(d2_71__N_490_adj_5690[24]), 
          .S1(d2_71__N_490_adj_5690[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_24 (.A0(d2_adj_5674[22]), .B0(d1_adj_5673[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[23]), .B1(d1_adj_5673[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15422), .COUT(n15423), .S0(d2_71__N_490_adj_5690[22]), 
          .S1(d2_71__N_490_adj_5690[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_22 (.A0(d2_adj_5674[20]), .B0(d1_adj_5673[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[21]), .B1(d1_adj_5673[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15421), .COUT(n15422), .S0(d2_71__N_490_adj_5690[20]), 
          .S1(d2_71__N_490_adj_5690[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_20 (.A0(d2_adj_5674[18]), .B0(d1_adj_5673[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[19]), .B1(d1_adj_5673[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15420), .COUT(n15421), .S0(d2_71__N_490_adj_5690[18]), 
          .S1(d2_71__N_490_adj_5690[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_18 (.A0(d2_adj_5674[16]), .B0(d1_adj_5673[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[17]), .B1(d1_adj_5673[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15419), .COUT(n15420), .S0(d2_71__N_490_adj_5690[16]), 
          .S1(d2_71__N_490_adj_5690[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_16 (.A0(d2_adj_5674[14]), .B0(d1_adj_5673[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[15]), .B1(d1_adj_5673[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15418), .COUT(n15419), .S0(d2_71__N_490_adj_5690[14]), 
          .S1(d2_71__N_490_adj_5690[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_14 (.A0(d2_adj_5674[12]), .B0(d1_adj_5673[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[13]), .B1(d1_adj_5673[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15417), .COUT(n15418), .S0(d2_71__N_490_adj_5690[12]), 
          .S1(d2_71__N_490_adj_5690[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_12 (.A0(d2_adj_5674[10]), .B0(d1_adj_5673[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[11]), .B1(d1_adj_5673[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15416), .COUT(n15417), .S0(d2_71__N_490_adj_5690[10]), 
          .S1(d2_71__N_490_adj_5690[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_10 (.A0(d2_adj_5674[8]), .B0(d1_adj_5673[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[9]), .B1(d1_adj_5673[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15415), .COUT(n15416), .S0(d2_71__N_490_adj_5690[8]), 
          .S1(d2_71__N_490_adj_5690[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_8 (.A0(d2_adj_5674[6]), .B0(d1_adj_5673[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[7]), .B1(d1_adj_5673[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15414), .COUT(n15415), .S0(d2_71__N_490_adj_5690[6]), 
          .S1(d2_71__N_490_adj_5690[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_6 (.A0(d2_adj_5674[4]), .B0(d1_adj_5673[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[5]), .B1(d1_adj_5673[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15413), .COUT(n15414), .S0(d2_71__N_490_adj_5690[4]), 
          .S1(d2_71__N_490_adj_5690[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_4 (.A0(d2_adj_5674[2]), .B0(d1_adj_5673[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[3]), .B1(d1_adj_5673[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15412), .COUT(n15413), .S0(d2_71__N_490_adj_5690[2]), 
          .S1(d2_71__N_490_adj_5690[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_2 (.A0(d2_adj_5674[0]), .B0(d1_adj_5673[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5674[1]), .B1(d1_adj_5673[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15412), .S1(d2_71__N_490_adj_5690[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1433_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_2.INJECT1_1 = "NO";
    LUT4 i5618_2_lut (.A(d2_adj_5674[0]), .B(d1_adj_5673[0]), .Z(d2_71__N_490_adj_5690[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5618_2_lut.init = 16'h6666;
    FD1S3AX phase_accum_e3_i0_i1 (.D(n318), .CK(clk_80mhz), .Q(phase_accum_adj_5665[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_1517_add_4_37 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n81_adj_5096), .D0(d1[70]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n78_adj_5095), .D1(d1[71]), .CIN(n15409), .S0(d1_71__N_418[70]), 
          .S1(d1_71__N_418[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_35 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n87_adj_5098), .D0(d1[68]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n84_adj_5097), .D1(d1[69]), .CIN(n15408), .COUT(n15409), 
          .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_33 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n93_adj_5100), .D0(d1[66]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n90_adj_5099), .D1(d1[67]), .CIN(n15407), .COUT(n15408), 
          .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_31 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n99_adj_5102), .D0(d1[64]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n96_adj_5101), .D1(d1[65]), .CIN(n15406), .COUT(n15407), 
          .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_29 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n105_adj_5104), .D0(d1[62]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n102_adj_5103), .D1(d1[63]), .CIN(n15405), .COUT(n15406), 
          .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_27 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n111_adj_5106), .D0(d1[60]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n108_adj_5105), .D1(d1[61]), .CIN(n15404), .COUT(n15405), 
          .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_25 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n117_adj_5108), .D0(d1[58]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n114_adj_5107), .D1(d1[59]), .CIN(n15403), .COUT(n15404), 
          .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_23 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n123_adj_5110), .D0(d1[56]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n120_adj_5109), .D1(d1[57]), .CIN(n15402), .COUT(n15403), 
          .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_21 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n129_adj_5112), .D0(d1[54]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n126_adj_5111), .D1(d1[55]), .CIN(n15401), .COUT(n15402), 
          .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_19 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n135_adj_5114), .D0(d1[52]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n132_adj_5113), .D1(d1[53]), .CIN(n15400), .COUT(n15401), 
          .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_11 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n159_adj_5122), .D0(d1[44]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n156_adj_5121), .D1(d1[45]), .CIN(n15396), .COUT(n15397), 
          .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_11.INJECT1_1 = "NO";
    LUT4 i5663_2_lut (.A(d3_adj_5675[0]), .B(d2_adj_5674[0]), .Z(d3_71__N_562_adj_5691[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5663_2_lut.init = 16'h6666;
    CCU2C _add_1_1517_add_4_17 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n141_adj_5116), .D0(d1[50]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n138_adj_5115), .D1(d1[51]), .CIN(n15399), .COUT(n15400), 
          .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_7 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n171_adj_5126), .D0(d1[40]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n168_adj_5125), .D1(d1[41]), .CIN(n15394), .COUT(n15395), 
          .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_15 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n147_adj_5118), .D0(d1[48]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n144_adj_5117), .D1(d1[49]), .CIN(n15398), .COUT(n15399), 
          .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_5 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n177_adj_5128), .D0(d1[38]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n174_adj_5127), .D1(d1[39]), .CIN(n15393), .COUT(n15394), 
          .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_3 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n183_adj_5130), .D0(d1[36]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n180_adj_5129), .D1(d1[37]), .CIN(n15392), .COUT(n15393), 
          .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_3.INJECT1_1 = "NO";
    LUT4 i2332_3_lut_4_lut (.A(n18138), .B(n18267), .C(led_c_3), .D(n154), 
         .Z(n12047)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2332_3_lut_4_lut.init = 16'hf707;
    CCU2C _add_1_1517_add_4_9 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n165_adj_5124), .D0(d1[42]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n162_adj_5123), .D1(d1[43]), .CIN(n15395), .COUT(n15396), 
          .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_13 (.A0(MixerOutSin[11]), .B0(cout_adj_5663), 
          .C0(n153_adj_5120), .D0(d1[46]), .A1(MixerOutSin[11]), .B1(cout_adj_5663), 
          .C1(n150_adj_5119), .D1(d1[47]), .CIN(n15397), .COUT(n15398), 
          .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_30 (.A0(d_d7[27]), .B0(d7[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[28]), .B1(d7[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16236), .COUT(n16237), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_30.INJECT1_1 = "NO";
    CCU2C add_4099_19 (.A0(d_out_d_11__N_1890[17]), .B0(n48_adj_5561), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n45_adj_5560), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16889), .S0(n912), .S1(d_out_d_11__N_1892[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_19.INIT0 = 16'h9995;
    defparam add_4099_19.INIT1 = 16'h9995;
    defparam add_4099_19.INJECT1_0 = "NO";
    defparam add_4099_19.INJECT1_1 = "NO";
    CCU2C add_4099_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1890[17]), .C0(n54_adj_5563), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n51_adj_5562), .D1(VCC_net), .CIN(n16888), .COUT(n16889), 
          .S0(n914), .S1(n913));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_17.INIT0 = 16'h6969;
    defparam add_4099_17.INIT1 = 16'h6969;
    defparam add_4099_17.INJECT1_0 = "NO";
    defparam add_4099_17.INJECT1_1 = "NO";
    CCU2C add_4099_15 (.A0(d_out_d_11__N_1890[17]), .B0(n60_adj_5565), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n57_adj_5564), .D1(VCC_net), .CIN(n16887), .COUT(n16888), 
          .S0(n916), .S1(n915));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_15.INIT0 = 16'h9995;
    defparam add_4099_15.INIT1 = 16'h6969;
    defparam add_4099_15.INJECT1_0 = "NO";
    defparam add_4099_15.INJECT1_1 = "NO";
    CCU2C add_4099_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n66_adj_5567), .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), 
          .B1(n18143), .C1(n63_adj_5566), .D1(VCC_net), .CIN(n16886), 
          .COUT(n16887), .S0(n918), .S1(n917));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_13.INIT0 = 16'h9696;
    defparam add_4099_13.INIT1 = 16'h6969;
    defparam add_4099_13.INJECT1_0 = "NO";
    defparam add_4099_13.INJECT1_1 = "NO";
    CCU2C add_4099_11 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n72_adj_5569), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n69_adj_5568), .D1(VCC_net), 
          .CIN(n16885), .COUT(n16886), .S0(n920), .S1(n919));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_11.INIT0 = 16'h9696;
    defparam add_4099_11.INIT1 = 16'h9696;
    defparam add_4099_11.INJECT1_0 = "NO";
    defparam add_4099_11.INJECT1_1 = "NO";
    CCU2C add_4099_9 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n78_adj_5571), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n75_adj_5570), .D1(VCC_net), 
          .CIN(n16884), .COUT(n16885), .S0(n922), .S1(n921));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_9.INIT0 = 16'h9696;
    defparam add_4099_9.INIT1 = 16'h9696;
    defparam add_4099_9.INJECT1_0 = "NO";
    defparam add_4099_9.INJECT1_1 = "NO";
    CCU2C add_4099_7 (.A0(d_out_d_11__N_1886[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n84_adj_5573), .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n81_adj_5572), .D1(VCC_net), 
          .CIN(n16883), .COUT(n16884), .S0(n924), .S1(n923));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_7.INIT0 = 16'h9696;
    defparam add_4099_7.INIT1 = 16'h9696;
    defparam add_4099_7.INJECT1_0 = "NO";
    defparam add_4099_7.INJECT1_1 = "NO";
    CCU2C add_4099_5 (.A0(n90_adj_5575), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(d_out_d_11__N_1890[17]), .C1(n87_adj_5574), 
          .D1(VCC_net), .CIN(n16882), .COUT(n16883), .S0(n926), .S1(n925));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_5.INIT0 = 16'haaa0;
    defparam add_4099_5.INIT1 = 16'h9696;
    defparam add_4099_5.INJECT1_0 = "NO";
    defparam add_4099_5.INJECT1_1 = "NO";
    CCU2C add_4099_3 (.A0(d_out_d_11__N_1890[17]), .B0(ISquare[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16881), .COUT(n16882), .S1(n927));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_3.INIT0 = 16'h666a;
    defparam add_4099_3.INIT1 = 16'h555f;
    defparam add_4099_3.INJECT1_0 = "NO";
    defparam add_4099_3.INJECT1_1 = "NO";
    CCU2C add_4099_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1890[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16881));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4099_1.INIT0 = 16'h0000;
    defparam add_4099_1.INIT1 = 16'haaaf;
    defparam add_4099_1.INJECT1_0 = "NO";
    defparam add_4099_1.INJECT1_1 = "NO";
    CCU2C add_4102_19 (.A0(d_out_d_11__N_1879), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1879), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16875), .S0(n45_adj_5513), 
          .S1(d_out_d_11__N_1882[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_19.INIT0 = 16'h666a;
    defparam add_4102_19.INIT1 = 16'h666a;
    defparam add_4102_19.INJECT1_0 = "NO";
    defparam add_4102_19.INJECT1_1 = "NO";
    CCU2C add_4102_17 (.A0(d_out_d_11__N_1880[17]), .B0(n54_adj_5305), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n51_adj_5304), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16874), .COUT(n16875), .S0(n51_adj_5515), 
          .S1(n48_adj_5514));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_17.INIT0 = 16'h9995;
    defparam add_4102_17.INIT1 = 16'h9995;
    defparam add_4102_17.INJECT1_0 = "NO";
    defparam add_4102_17.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_28 (.A0(d_d7[25]), .B0(d7[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[26]), .B1(d7[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16235), .COUT(n16236), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_28.INJECT1_1 = "NO";
    CCU2C add_4102_15 (.A0(d_out_d_11__N_1880[17]), .B0(n60_adj_5307), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n57_adj_5306), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16873), .COUT(n16874), .S0(n57_adj_5517), 
          .S1(n54_adj_5516));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_15.INIT0 = 16'h9995;
    defparam add_4102_15.INIT1 = 16'h9995;
    defparam add_4102_15.INJECT1_0 = "NO";
    defparam add_4102_15.INJECT1_1 = "NO";
    CCU2C add_4102_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n66_adj_5309), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n63_adj_5308), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16872), .COUT(n16873), .S0(n63_adj_5519), 
          .S1(n60_adj_5518));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_13.INIT0 = 16'h6969;
    defparam add_4102_13.INIT1 = 16'h9995;
    defparam add_4102_13.INJECT1_0 = "NO";
    defparam add_4102_13.INJECT1_1 = "NO";
    CCU2C add_4102_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n72_adj_5311), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1880[17]), 
          .C1(n69_adj_5310), .D1(VCC_net), .CIN(n16871), .COUT(n16872), 
          .S0(n69_adj_5521), .S1(n66_adj_5520));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_11.INIT0 = 16'h6969;
    defparam add_4102_11.INIT1 = 16'h6969;
    defparam add_4102_11.INJECT1_0 = "NO";
    defparam add_4102_11.INJECT1_1 = "NO";
    CCU2C add_4102_9 (.A0(d_out_d_11__N_1880[17]), .B0(n18143), .C0(n78_adj_5313), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n75_adj_5312), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16870), .COUT(n16871), .S0(n75_adj_5523), 
          .S1(n72_adj_5522));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_9.INIT0 = 16'h6969;
    defparam add_4102_9.INIT1 = 16'h9995;
    defparam add_4102_9.INJECT1_0 = "NO";
    defparam add_4102_9.INJECT1_1 = "NO";
    CCU2C add_4102_7 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(n84_adj_5315), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1880[17]), .C1(n81_adj_5314), .D1(VCC_net), 
          .CIN(n16869), .COUT(n16870), .S0(n81_adj_5525), .S1(n78_adj_5524));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_7.INIT0 = 16'h9696;
    defparam add_4102_7.INIT1 = 16'h9696;
    defparam add_4102_7.INJECT1_0 = "NO";
    defparam add_4102_7.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_18 (.A0(d4_adj_5676[51]), .B0(d3_adj_5675[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[52]), .B1(d3_adj_5675[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16275), .COUT(n16276), .S0(n138_adj_4741), 
          .S1(n135_adj_4791));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_18.INJECT1_1 = "NO";
    CCU2C add_4102_5 (.A0(n90_adj_5317), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1880[17]), .C1(n87_adj_5316), 
          .D1(VCC_net), .CIN(n16868), .COUT(n16869), .S0(n87_adj_5527), 
          .S1(n84_adj_5526));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_5.INIT0 = 16'haaa0;
    defparam add_4102_5.INIT1 = 16'h9696;
    defparam add_4102_5.INJECT1_0 = "NO";
    defparam add_4102_5.INJECT1_1 = "NO";
    CCU2C add_4102_3 (.A0(d_out_d_11__N_1880[17]), .B0(ISquare[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16867), .COUT(n16868), .S1(n90_adj_5528));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_3.INIT0 = 16'h666a;
    defparam add_4102_3.INIT1 = 16'h555f;
    defparam add_4102_3.INJECT1_0 = "NO";
    defparam add_4102_3.INJECT1_1 = "NO";
    CCU2C add_4102_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16867));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4102_1.INIT0 = 16'h0000;
    defparam add_4102_1.INIT1 = 16'haaaf;
    defparam add_4102_1.INJECT1_0 = "NO";
    defparam add_4102_1.INJECT1_1 = "NO";
    CCU2C add_4103_19 (.A0(d_out_d_11__N_1884[17]), .B0(n48_adj_5530), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n45_adj_5529), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16861), .S0(n45_adj_5497), 
          .S1(d_out_d_11__N_1886[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_19.INIT0 = 16'h9995;
    defparam add_4103_19.INIT1 = 16'h9995;
    defparam add_4103_19.INJECT1_0 = "NO";
    defparam add_4103_19.INJECT1_1 = "NO";
    LUT4 i6627_4_lut (.A(n18301), .B(led_c_3), .C(n13099), .D(n18141), 
         .Z(clk_80mhz_enable_1471)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;
    defparam i6627_4_lut.init = 16'ha0a2;
    CCU2C add_4103_17 (.A0(d_out_d_11__N_1884[17]), .B0(n54_adj_5532), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n51_adj_5531), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16860), .COUT(n16861), .S0(n51_adj_5499), 
          .S1(n48_adj_5498));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_17.INIT0 = 16'h9995;
    defparam add_4103_17.INIT1 = 16'h9995;
    defparam add_4103_17.INJECT1_0 = "NO";
    defparam add_4103_17.INJECT1_1 = "NO";
    CCU2C add_4103_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n60_adj_5534), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n57_adj_5533), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16859), .COUT(n16860), .S0(n57_adj_5501), 
          .S1(n54_adj_5500));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_15.INIT0 = 16'h6969;
    defparam add_4103_15.INIT1 = 16'h9995;
    defparam add_4103_15.INJECT1_0 = "NO";
    defparam add_4103_15.INJECT1_1 = "NO";
    CCU2C add_4103_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n66_adj_5536), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1884[17]), 
          .C1(n63_adj_5535), .D1(VCC_net), .CIN(n16858), .COUT(n16859), 
          .S0(n63_adj_5503), .S1(n60_adj_5502));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_13.INIT0 = 16'h6969;
    defparam add_4103_13.INIT1 = 16'h6969;
    defparam add_4103_13.INJECT1_0 = "NO";
    defparam add_4103_13.INJECT1_1 = "NO";
    CCU2C add_4103_11 (.A0(d_out_d_11__N_1884[17]), .B0(n18143), .C0(n72_adj_5538), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n69_adj_5537), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16857), .COUT(n16858), .S0(n69_adj_5505), 
          .S1(n66_adj_5504));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_11.INIT0 = 16'h6969;
    defparam add_4103_11.INIT1 = 16'h9995;
    defparam add_4103_11.INJECT1_0 = "NO";
    defparam add_4103_11.INJECT1_1 = "NO";
    CCU2C add_4103_9 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n78_adj_5540), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n75_adj_5539), .D1(VCC_net), 
          .CIN(n16856), .COUT(n16857), .S0(n75_adj_5507), .S1(n72_adj_5506));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_9.INIT0 = 16'h9696;
    defparam add_4103_9.INIT1 = 16'h9696;
    defparam add_4103_9.INJECT1_0 = "NO";
    defparam add_4103_9.INJECT1_1 = "NO";
    CCU2C add_4103_7 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n84_adj_5542), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n81_adj_5541), .D1(VCC_net), 
          .CIN(n16855), .COUT(n16856), .S0(n81_adj_5509), .S1(n78_adj_5508));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_7.INIT0 = 16'h9696;
    defparam add_4103_7.INIT1 = 16'h9696;
    defparam add_4103_7.INJECT1_0 = "NO";
    defparam add_4103_7.INJECT1_1 = "NO";
    CCU2C add_4103_5 (.A0(n90_adj_5544), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(d_out_d_11__N_1884[17]), .C1(n87_adj_5543), 
          .D1(VCC_net), .CIN(n16854), .COUT(n16855), .S0(n87_adj_5511), 
          .S1(n84_adj_5510));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_5.INIT0 = 16'haaa0;
    defparam add_4103_5.INIT1 = 16'h9696;
    defparam add_4103_5.INJECT1_0 = "NO";
    defparam add_4103_5.INJECT1_1 = "NO";
    CCU2C add_4103_3 (.A0(d_out_d_11__N_1884[17]), .B0(ISquare[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16853), .COUT(n16854), .S1(n90_adj_5512));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_3.INIT0 = 16'h666a;
    defparam add_4103_3.INIT1 = 16'h555f;
    defparam add_4103_3.INJECT1_0 = "NO";
    defparam add_4103_3.INJECT1_1 = "NO";
    CCU2C add_4103_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16853));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4103_1.INIT0 = 16'h0000;
    defparam add_4103_1.INIT1 = 16'haaaf;
    defparam add_4103_1.INJECT1_0 = "NO";
    defparam add_4103_1.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i2 (.D(n315), .CK(clk_80mhz), .Q(phase_accum_adj_5665[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i3 (.D(n312), .CK(clk_80mhz), .Q(phase_accum_adj_5665[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i4 (.D(n309), .CK(clk_80mhz), .Q(phase_accum_adj_5665[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i5 (.D(n306), .CK(clk_80mhz), .Q(phase_accum_adj_5665[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i6 (.D(n303), .CK(clk_80mhz), .Q(phase_accum_adj_5665[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i7 (.D(n300), .CK(clk_80mhz), .Q(phase_accum_adj_5665[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i8 (.D(n297), .CK(clk_80mhz), .Q(phase_accum_adj_5665[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i9 (.D(n294), .CK(clk_80mhz), .Q(phase_accum_adj_5665[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i10 (.D(n291), .CK(clk_80mhz), .Q(phase_accum_adj_5665[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i11 (.D(n288), .CK(clk_80mhz), .Q(phase_accum_adj_5665[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i12 (.D(n285), .CK(clk_80mhz), .Q(phase_accum_adj_5665[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i13 (.D(n282), .CK(clk_80mhz), .Q(phase_accum_adj_5665[13]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i14 (.D(n279), .CK(clk_80mhz), .Q(phase_accum_adj_5665[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i15 (.D(n276), .CK(clk_80mhz), .Q(phase_accum_adj_5665[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i16 (.D(n273), .CK(clk_80mhz), .Q(phase_accum_adj_5665[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i17 (.D(n270), .CK(clk_80mhz), .Q(phase_accum_adj_5665[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i18 (.D(n267), .CK(clk_80mhz), .Q(phase_accum_adj_5665[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i19 (.D(n264), .CK(clk_80mhz), .Q(phase_accum_adj_5665[19]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i20 (.D(n261), .CK(clk_80mhz), .Q(phase_accum_adj_5665[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i21 (.D(n258), .CK(clk_80mhz), .Q(phase_accum_adj_5665[21]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i22 (.D(n255), .CK(clk_80mhz), .Q(phase_accum_adj_5665[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i23 (.D(n252), .CK(clk_80mhz), .Q(phase_accum_adj_5665[23]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i24 (.D(n249), .CK(clk_80mhz), .Q(phase_accum_adj_5665[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i25 (.D(n246), .CK(clk_80mhz), .Q(phase_accum_adj_5665[25]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i26 (.D(n243), .CK(clk_80mhz), .Q(phase_accum_adj_5665[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i27 (.D(n240), .CK(clk_80mhz), .Q(phase_accum_adj_5665[27]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i28 (.D(n237), .CK(clk_80mhz), .Q(phase_accum_adj_5665[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i29 (.D(n234), .CK(clk_80mhz), .Q(phase_accum_adj_5665[29]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i30 (.D(n231), .CK(clk_80mhz), .Q(phase_accum_adj_5665[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i31 (.D(n228), .CK(clk_80mhz), .Q(phase_accum_adj_5665[31]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i32 (.D(n225), .CK(clk_80mhz), .Q(phase_accum_adj_5665[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i33 (.D(n222), .CK(clk_80mhz), .Q(phase_accum_adj_5665[33]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i34 (.D(n219), .CK(clk_80mhz), .Q(phase_accum_adj_5665[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i35 (.D(n216), .CK(clk_80mhz), .Q(phase_accum_adj_5665[35]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i36 (.D(n213), .CK(clk_80mhz), .Q(phase_accum_adj_5665[36]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i37 (.D(n210), .CK(clk_80mhz), .Q(phase_accum_adj_5665[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i38 (.D(n207), .CK(clk_80mhz), .Q(phase_accum_adj_5665[38]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i39 (.D(n204), .CK(clk_80mhz), .Q(phase_accum_adj_5665[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i40 (.D(n201), .CK(clk_80mhz), .Q(phase_accum_adj_5665[40]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i41 (.D(n198), .CK(clk_80mhz), .Q(phase_accum_adj_5665[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i42 (.D(n195), .CK(clk_80mhz), .Q(phase_accum_adj_5665[42]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i43 (.D(n192), .CK(clk_80mhz), .Q(phase_accum_adj_5665[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i44 (.D(n189), .CK(clk_80mhz), .Q(phase_accum_adj_5665[44]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i45 (.D(n186), .CK(clk_80mhz), .Q(phase_accum_adj_5665[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i46 (.D(n183_adj_4733), .CK(clk_80mhz), .Q(phase_accum_adj_5665[46]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i47 (.D(n180_adj_4734), .CK(clk_80mhz), .Q(phase_accum_adj_5665[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i48 (.D(n177_adj_4735), .CK(clk_80mhz), .Q(phase_accum_adj_5665[48]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i49 (.D(n174_adj_4737), .CK(clk_80mhz), .Q(phase_accum_adj_5665[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i50 (.D(n171_adj_4738), .CK(clk_80mhz), .Q(phase_accum_adj_5665[50]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i51 (.D(n168_adj_4743), .CK(clk_80mhz), .Q(phase_accum_adj_5665[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i52 (.D(n165_adj_4748), .CK(clk_80mhz), .Q(phase_accum_adj_5665[52]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i53 (.D(n162_adj_4749), .CK(clk_80mhz), .Q(phase_accum_adj_5665[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i54 (.D(n159_adj_4750), .CK(clk_80mhz), .Q(phase_accum_adj_5665[54]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i55 (.D(n156_adj_4751), .CK(clk_80mhz), .Q(phase_accum_adj_5665[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i56 (.D(n153_adj_4752), .CK(clk_80mhz), .Q(phase_accum[56]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i57 (.D(n150_adj_4753), .CK(clk_80mhz), .Q(phase_accum[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i58 (.D(n147_adj_4754), .CK(clk_80mhz), .Q(phase_accum[58]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i59 (.D(n144_adj_4769), .CK(clk_80mhz), .Q(phase_accum[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i60 (.D(n141_adj_4784), .CK(clk_80mhz), .Q(phase_accum[60]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i61 (.D(n138_adj_4785), .CK(clk_80mhz), .Q(phase_accum[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i62 (.D(n135_adj_4786), .CK(clk_80mhz), .Q(phase_accum[62]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i63 (.D(n132_adj_4787), .CK(clk_80mhz), .Q(phase_accum[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_1628_add_4_4 (.A0(d_d6_adj_5679[37]), .B0(d6_adj_5678[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5679[38]), .B1(d6_adj_5678[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16664), .COUT(n16665), .S0(n180_adj_5388), 
          .S1(n177_adj_5387));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_4.INJECT1_1 = "NO";
    CCU2C add_4104_17 (.A0(d_out_d_11__N_1877), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1877), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16847), .S0(n51_adj_5304), 
          .S1(d_out_d_11__N_1880[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_17.INIT0 = 16'h666a;
    defparam add_4104_17.INIT1 = 16'h666a;
    defparam add_4104_17.INJECT1_0 = "NO";
    defparam add_4104_17.INJECT1_1 = "NO";
    CCU2C add_4104_15 (.A0(d_out_d_11__N_1878[17]), .B0(n55), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n52), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16846), .COUT(n16847), .S0(n57_adj_5306), 
          .S1(n54_adj_5305));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_15.INIT0 = 16'h9995;
    defparam add_4104_15.INIT1 = 16'h9995;
    defparam add_4104_15.INJECT1_0 = "NO";
    defparam add_4104_15.INJECT1_1 = "NO";
    CCU2C add_4104_13 (.A0(d_out_d_11__N_1878[17]), .B0(n61), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n58), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16845), .COUT(n16846), .S0(n63_adj_5308), 
          .S1(n60_adj_5307));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_13.INIT0 = 16'h9995;
    defparam add_4104_13.INIT1 = 16'h9995;
    defparam add_4104_13.INJECT1_0 = "NO";
    defparam add_4104_13.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5679[36]), .B1(d6_adj_5678[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16664), .S1(n183_adj_5389));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1628_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1628_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_2.INJECT1_1 = "NO";
    CCU2C add_4104_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1878[17]), .C0(n67), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n64_adj_5491), .D1(VCC_net), .CIN(n16844), .COUT(n16845), 
          .S0(n69_adj_5310), .S1(n66_adj_5309));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_11.INIT0 = 16'h6969;
    defparam add_4104_11.INIT1 = 16'h6969;
    defparam add_4104_11.INJECT1_0 = "NO";
    defparam add_4104_11.INJECT1_1 = "NO";
    CCU2C add_4104_9 (.A0(d_out_d_11__N_1878[17]), .B0(n73), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n70), .D1(VCC_net), .CIN(n16843), .COUT(n16844), .S0(n75_adj_5312), 
          .S1(n72_adj_5311));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_9.INIT0 = 16'h9995;
    defparam add_4104_9.INIT1 = 16'h6969;
    defparam add_4104_9.INJECT1_0 = "NO";
    defparam add_4104_9.INJECT1_1 = "NO";
    CCU2C add_4104_7 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1878[17]), 
          .C0(n79_adj_5493), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(n18143), .C1(n76_adj_5492), .D1(VCC_net), .CIN(n16842), 
          .COUT(n16843), .S0(n81_adj_5314), .S1(n78_adj_5313));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_7.INIT0 = 16'h9696;
    defparam add_4104_7.INIT1 = 16'h6969;
    defparam add_4104_7.INJECT1_0 = "NO";
    defparam add_4104_7.INJECT1_1 = "NO";
    CCU2C add_4104_5 (.A0(n85_adj_5495), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1878[17]), .C1(n82_adj_5494), 
          .D1(VCC_net), .CIN(n16841), .COUT(n16842), .S0(n87_adj_5316), 
          .S1(n84_adj_5315));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_5.INIT0 = 16'haaa0;
    defparam add_4104_5.INIT1 = 16'h9696;
    defparam add_4104_5.INJECT1_0 = "NO";
    defparam add_4104_5.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_63 (.A0(phase_inc_carrGen[62]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16662), .S0(n133_adj_5391), 
          .S1(n130_adj_5390));
    defparam _add_1_1457_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_63.INJECT1_1 = "NO";
    CCU2C add_4104_3 (.A0(d_out_d_11__N_1878[17]), .B0(ISquare[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16840), .COUT(n16841), .S1(n90_adj_5317));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_3.INIT0 = 16'h666a;
    defparam add_4104_3.INIT1 = 16'h555f;
    defparam add_4104_3.INJECT1_0 = "NO";
    defparam add_4104_3.INJECT1_1 = "NO";
    CCU2C add_4104_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16840));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4104_1.INIT0 = 16'h0000;
    defparam add_4104_1.INIT1 = 16'haaaf;
    defparam add_4104_1.INJECT1_0 = "NO";
    defparam add_4104_1.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_61 (.A0(phase_inc_carrGen[60]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16661), .COUT(n16662), .S0(n139_adj_5393), 
          .S1(n136_adj_5392));
    defparam _add_1_1457_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_61.INJECT1_1 = "NO";
    CCU2C add_4108_15 (.A0(d_out_d_11__N_1875), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1875), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16834), .S0(n52), .S1(d_out_d_11__N_1878[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_15.INIT0 = 16'h666a;
    defparam add_4108_15.INIT1 = 16'h666a;
    defparam add_4108_15.INJECT1_0 = "NO";
    defparam add_4108_15.INJECT1_1 = "NO";
    CCU2C add_4108_13 (.A0(d_out_d_11__N_1876[17]), .B0(n51_adj_5614), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n48_adj_5613), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16833), .COUT(n16834), .S0(n58), 
          .S1(n55));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_13.INIT0 = 16'h9995;
    defparam add_4108_13.INIT1 = 16'h9995;
    defparam add_4108_13.INJECT1_0 = "NO";
    defparam add_4108_13.INJECT1_1 = "NO";
    CCU2C add_4108_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n57_adj_5616), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n54_adj_5615), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16832), .COUT(n16833), .S0(n64_adj_5491), 
          .S1(n61));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_11.INIT0 = 16'h6969;
    defparam add_4108_11.INIT1 = 16'h9995;
    defparam add_4108_11.INJECT1_0 = "NO";
    defparam add_4108_11.INJECT1_1 = "NO";
    CCU2C add_4108_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n63_adj_5618), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1876[17]), 
          .C1(n60_adj_5617), .D1(VCC_net), .CIN(n16831), .COUT(n16832), 
          .S0(n70), .S1(n67));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_9.INIT0 = 16'h6969;
    defparam add_4108_9.INIT1 = 16'h6969;
    defparam add_4108_9.INJECT1_0 = "NO";
    defparam add_4108_9.INJECT1_1 = "NO";
    CCU2C add_4108_7 (.A0(d_out_d_11__N_1876[17]), .B0(n18143), .C0(n69_adj_5620), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n66_adj_5619), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16830), .COUT(n16831), .S0(n76_adj_5492), 
          .S1(n73));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_7.INIT0 = 16'h6969;
    defparam add_4108_7.INIT1 = 16'h9995;
    defparam add_4108_7.INJECT1_0 = "NO";
    defparam add_4108_7.INJECT1_1 = "NO";
    CCU2C add_4108_5 (.A0(n75_adj_5622), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1876[17]), .C1(n72_adj_5621), 
          .D1(VCC_net), .CIN(n16829), .COUT(n16830), .S0(n82_adj_5494), 
          .S1(n79_adj_5493));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_5.INIT0 = 16'haaa0;
    defparam add_4108_5.INIT1 = 16'h9696;
    defparam add_4108_5.INJECT1_0 = "NO";
    defparam add_4108_5.INJECT1_1 = "NO";
    CCU2C add_4108_3 (.A0(d_out_d_11__N_1876[17]), .B0(ISquare[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16828), .COUT(n16829), .S1(n85_adj_5495));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_3.INIT0 = 16'h666a;
    defparam add_4108_3.INIT1 = 16'h555f;
    defparam add_4108_3.INJECT1_0 = "NO";
    defparam add_4108_3.INJECT1_1 = "NO";
    CCU2C add_4108_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16828));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4108_1.INIT0 = 16'h0000;
    defparam add_4108_1.INIT1 = 16'haaaf;
    defparam add_4108_1.INJECT1_0 = "NO";
    defparam add_4108_1.INJECT1_1 = "NO";
    CCU2C add_4109_17 (.A0(ISquare[31]), .B0(n913), .C0(GND_net), .D0(VCC_net), 
          .A1(n912), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16822), 
          .S1(d_out_d_11__N_2353[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_17.INIT0 = 16'h666a;
    defparam add_4109_17.INIT1 = 16'haaa0;
    defparam add_4109_17.INJECT1_0 = "NO";
    defparam add_4109_17.INJECT1_1 = "NO";
    CCU2C add_4109_15 (.A0(ISquare[31]), .B0(n915), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n914), .C1(GND_net), .D1(VCC_net), .CIN(n16821), 
          .COUT(n16822));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_15.INIT0 = 16'h666a;
    defparam add_4109_15.INIT1 = 16'h666a;
    defparam add_4109_15.INJECT1_0 = "NO";
    defparam add_4109_15.INJECT1_1 = "NO";
    CCU2C add_4109_13 (.A0(n917), .B0(n15364), .C0(n209), .D0(ISquare[31]), 
          .A1(n916), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16820), 
          .COUT(n16821));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_13.INIT0 = 16'h556a;
    defparam add_4109_13.INIT1 = 16'haaa0;
    defparam add_4109_13.INJECT1_0 = "NO";
    defparam add_4109_13.INJECT1_1 = "NO";
    CCU2C add_4109_11 (.A0(d_out_d_11__N_1876[17]), .B0(n919), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n918), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16819), .COUT(n16820));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_11.INIT0 = 16'h9995;
    defparam add_4109_11.INIT1 = 16'h9995;
    defparam add_4109_11.INJECT1_0 = "NO";
    defparam add_4109_11.INJECT1_1 = "NO";
    CCU2C add_4109_9 (.A0(d_out_d_11__N_1880[17]), .B0(n921), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n920), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16818), .COUT(n16819));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_9.INIT0 = 16'h9995;
    defparam add_4109_9.INIT1 = 16'h9995;
    defparam add_4109_9.INJECT1_0 = "NO";
    defparam add_4109_9.INJECT1_1 = "NO";
    CCU2C add_4109_7 (.A0(d_out_d_11__N_1884[17]), .B0(n923), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n922), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16817), .COUT(n16818));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_7.INIT0 = 16'h9995;
    defparam add_4109_7.INIT1 = 16'h9995;
    defparam add_4109_7.INJECT1_0 = "NO";
    defparam add_4109_7.INJECT1_1 = "NO";
    CCU2C add_4109_5 (.A0(d_out_d_11__N_1888[17]), .B0(n925), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n924), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16816), .COUT(n16817));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_5.INIT0 = 16'h9995;
    defparam add_4109_5.INIT1 = 16'h9995;
    defparam add_4109_5.INJECT1_0 = "NO";
    defparam add_4109_5.INJECT1_1 = "NO";
    CCU2C add_4109_3 (.A0(d_out_d_11__N_1892[17]), .B0(n927), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n926), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16815), .COUT(n16816));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_3.INIT0 = 16'h9995;
    defparam add_4109_3.INIT1 = 16'h9995;
    defparam add_4109_3.INJECT1_0 = "NO";
    defparam add_4109_3.INJECT1_1 = "NO";
    CCU2C add_4109_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(ISquare[0]), 
          .A1(d_out_d_11__N_1892[17]), .B1(ISquare[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16815));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(58[15:27])
    defparam add_4109_1.INIT0 = 16'h000A;
    defparam add_4109_1.INIT1 = 16'h666a;
    defparam add_4109_1.INJECT1_0 = "NO";
    defparam add_4109_1.INJECT1_1 = "NO";
    CCU2C add_4100_19 (.A0(d_out_d_11__N_1882[17]), .B0(n48_adj_5514), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n45_adj_5513), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16813), .S0(n45_adj_5529), 
          .S1(d_out_d_11__N_1884[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_19.INIT0 = 16'h9995;
    defparam add_4100_19.INIT1 = 16'h9995;
    defparam add_4100_19.INJECT1_0 = "NO";
    defparam add_4100_19.INJECT1_1 = "NO";
    CCU2C add_4100_17 (.A0(d_out_d_11__N_1882[17]), .B0(n54_adj_5516), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n51_adj_5515), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16812), .COUT(n16813), .S0(n51_adj_5531), 
          .S1(n48_adj_5530));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_17.INIT0 = 16'h9995;
    defparam add_4100_17.INIT1 = 16'h9995;
    defparam add_4100_17.INJECT1_0 = "NO";
    defparam add_4100_17.INJECT1_1 = "NO";
    CCU2C add_4100_15 (.A0(d_out_d_11__N_1882[17]), .B0(n60_adj_5518), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n57_adj_5517), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16811), .COUT(n16812), .S0(n57_adj_5533), 
          .S1(n54_adj_5532));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_15.INIT0 = 16'h9995;
    defparam add_4100_15.INIT1 = 16'h9995;
    defparam add_4100_15.INJECT1_0 = "NO";
    defparam add_4100_15.INJECT1_1 = "NO";
    CCU2C add_4100_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1882[17]), .C0(n66_adj_5520), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n63_adj_5519), .D1(VCC_net), .CIN(n16810), .COUT(n16811), 
          .S0(n63_adj_5535), .S1(n60_adj_5534));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_13.INIT0 = 16'h6969;
    defparam add_4100_13.INIT1 = 16'h6969;
    defparam add_4100_13.INJECT1_0 = "NO";
    defparam add_4100_13.INJECT1_1 = "NO";
    CCU2C add_4100_11 (.A0(d_out_d_11__N_1882[17]), .B0(n72_adj_5522), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n69_adj_5521), .D1(VCC_net), .CIN(n16809), .COUT(n16810), 
          .S0(n69_adj_5537), .S1(n66_adj_5536));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_11.INIT0 = 16'h9995;
    defparam add_4100_11.INIT1 = 16'h6969;
    defparam add_4100_11.INJECT1_0 = "NO";
    defparam add_4100_11.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_59 (.A0(phase_inc_carrGen[58]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16660), .COUT(n16661), .S0(n145_adj_5395), 
          .S1(n142_adj_5394));
    defparam _add_1_1457_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_59.INJECT1_1 = "NO";
    CCU2C add_4100_9 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n78_adj_5524), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(n18143), .C1(n75_adj_5523), .D1(VCC_net), .CIN(n16808), 
          .COUT(n16809), .S0(n75_adj_5539), .S1(n72_adj_5538));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_9.INIT0 = 16'h9696;
    defparam add_4100_9.INIT1 = 16'h6969;
    defparam add_4100_9.INJECT1_0 = "NO";
    defparam add_4100_9.INJECT1_1 = "NO";
    CCU2C add_4100_7 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n84_adj_5526), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(n81_adj_5525), .D1(VCC_net), 
          .CIN(n16807), .COUT(n16808), .S0(n81_adj_5541), .S1(n78_adj_5540));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_7.INIT0 = 16'h9696;
    defparam add_4100_7.INIT1 = 16'h9696;
    defparam add_4100_7.INJECT1_0 = "NO";
    defparam add_4100_7.INJECT1_1 = "NO";
    CCU2C add_4100_5 (.A0(n90_adj_5528), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1882[17]), .C1(n87_adj_5527), 
          .D1(VCC_net), .CIN(n16806), .COUT(n16807), .S0(n87_adj_5543), 
          .S1(n84_adj_5542));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_5.INIT0 = 16'haaa0;
    defparam add_4100_5.INIT1 = 16'h9696;
    defparam add_4100_5.INJECT1_0 = "NO";
    defparam add_4100_5.INJECT1_1 = "NO";
    CCU2C add_4100_3 (.A0(d_out_d_11__N_1882[17]), .B0(ISquare[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16805), .COUT(n16806), .S1(n90_adj_5544));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_3.INIT0 = 16'h666a;
    defparam add_4100_3.INIT1 = 16'h555f;
    defparam add_4100_3.INJECT1_0 = "NO";
    defparam add_4100_3.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_57 (.A0(phase_inc_carrGen[56]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16659), .COUT(n16660), .S0(n151_adj_5397), 
          .S1(n148_adj_5396));
    defparam _add_1_1457_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_57.INJECT1_1 = "NO";
    CCU2C add_4100_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16805));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4100_1.INIT0 = 16'h0000;
    defparam add_4100_1.INIT1 = 16'haaaf;
    defparam add_4100_1.INJECT1_0 = "NO";
    defparam add_4100_1.INJECT1_1 = "NO";
    CCU2C add_4110_19 (.A0(d_out_d_11__N_1886[17]), .B0(n48_adj_5498), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n45_adj_5497), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16799), .S0(n45_adj_5133), 
          .S1(d_out_d_11__N_1888[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_19.INIT0 = 16'h9995;
    defparam add_4110_19.INIT1 = 16'h9995;
    defparam add_4110_19.INJECT1_0 = "NO";
    defparam add_4110_19.INJECT1_1 = "NO";
    CCU2C add_4110_17 (.A0(d_out_d_11__N_1886[17]), .B0(n54_adj_5500), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n51_adj_5499), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16798), .COUT(n16799), .S0(n51_adj_5135), 
          .S1(n48_adj_5134));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_17.INIT0 = 16'h9995;
    defparam add_4110_17.INIT1 = 16'h9995;
    defparam add_4110_17.INJECT1_0 = "NO";
    defparam add_4110_17.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_55 (.A0(phase_inc_carrGen[54]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16658), .COUT(n16659), .S0(n157_adj_5399), 
          .S1(n154_adj_5398));
    defparam _add_1_1457_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_55.INJECT1_1 = "NO";
    CCU2C add_4110_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1886[17]), .C0(n60_adj_5502), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n57_adj_5501), .D1(VCC_net), .CIN(n16797), .COUT(n16798), 
          .S0(n57_adj_5137), .S1(n54_adj_5136));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_15.INIT0 = 16'h6969;
    defparam add_4110_15.INIT1 = 16'h6969;
    defparam add_4110_15.INJECT1_0 = "NO";
    defparam add_4110_15.INJECT1_1 = "NO";
    CCU2C add_4110_13 (.A0(d_out_d_11__N_1886[17]), .B0(n66_adj_5504), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n63_adj_5503), .D1(VCC_net), .CIN(n16796), .COUT(n16797), 
          .S0(n63_adj_5139), .S1(n60_adj_5138));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_13.INIT0 = 16'h9995;
    defparam add_4110_13.INIT1 = 16'h6969;
    defparam add_4110_13.INJECT1_0 = "NO";
    defparam add_4110_13.INJECT1_1 = "NO";
    CCU2C add_4110_11 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n72_adj_5506), .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), 
          .B1(n18143), .C1(n69_adj_5505), .D1(VCC_net), .CIN(n16795), 
          .COUT(n16796), .S0(n69_adj_5141), .S1(n66_adj_5140));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_11.INIT0 = 16'h9696;
    defparam add_4110_11.INIT1 = 16'h6969;
    defparam add_4110_11.INJECT1_0 = "NO";
    defparam add_4110_11.INJECT1_1 = "NO";
    CCU2C add_4110_9 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n78_adj_5508), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n75_adj_5507), .D1(VCC_net), 
          .CIN(n16794), .COUT(n16795), .S0(n75_adj_5143), .S1(n72_adj_5142));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_9.INIT0 = 16'h9696;
    defparam add_4110_9.INIT1 = 16'h9696;
    defparam add_4110_9.INJECT1_0 = "NO";
    defparam add_4110_9.INJECT1_1 = "NO";
    CCU2C add_4110_7 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n84_adj_5510), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n81_adj_5509), .D1(VCC_net), 
          .CIN(n16793), .COUT(n16794), .S0(n81_adj_5145), .S1(n78_adj_5144));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_7.INIT0 = 16'h9696;
    defparam add_4110_7.INIT1 = 16'h9696;
    defparam add_4110_7.INJECT1_0 = "NO";
    defparam add_4110_7.INJECT1_1 = "NO";
    CCU2C add_4110_5 (.A0(n90_adj_5512), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(d_out_d_11__N_1886[17]), .C1(n87_adj_5511), 
          .D1(VCC_net), .CIN(n16792), .COUT(n16793), .S0(n87_adj_5147), 
          .S1(n84_adj_5146));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_5.INIT0 = 16'haaa0;
    defparam add_4110_5.INIT1 = 16'h9696;
    defparam add_4110_5.INJECT1_0 = "NO";
    defparam add_4110_5.INJECT1_1 = "NO";
    CCU2C add_4110_3 (.A0(d_out_d_11__N_1886[17]), .B0(ISquare[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16791), .COUT(n16792), .S1(n90_adj_5148));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_3.INIT0 = 16'h666a;
    defparam add_4110_3.INIT1 = 16'h555f;
    defparam add_4110_3.INJECT1_0 = "NO";
    defparam add_4110_3.INJECT1_1 = "NO";
    CCU2C add_4110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16791));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4110_1.INIT0 = 16'h0000;
    defparam add_4110_1.INIT1 = 16'haaaf;
    defparam add_4110_1.INJECT1_0 = "NO";
    defparam add_4110_1.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_26 (.A0(d_d7[23]), .B0(d7[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[24]), .B1(d7[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16234), .COUT(n16235), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_24 (.A0(d_d7[21]), .B0(d7[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[22]), .B1(d7[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16233), .COUT(n16234), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_22 (.A0(d_d7[19]), .B0(d7[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[20]), .B1(d7[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16232), .COUT(n16233), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_20 (.A0(d_d7[17]), .B0(d7[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[18]), .B1(d7[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16231), .COUT(n16232), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_18 (.A0(d_d7[15]), .B0(d7[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[16]), .B1(d7[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16230), .COUT(n16231), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_16 (.A0(d_d7[13]), .B0(d7[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[14]), .B1(d7[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16229), .COUT(n16230), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_14 (.A0(d_d7[11]), .B0(d7[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[12]), .B1(d7[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16228), .COUT(n16229), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_12 (.A0(d_d7[9]), .B0(d7[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[10]), .B1(d7[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16227), .COUT(n16228), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_10 (.A0(d_d7[7]), .B0(d7[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[8]), .B1(d7[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16226), .COUT(n16227), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_8 (.A0(d_d7[5]), .B0(d7[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[6]), .B1(d7[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16225), .COUT(n16226), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_6 (.A0(d_d7[3]), .B0(d7[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[4]), .B1(d7[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16224), .COUT(n16225), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_4 (.A0(d_d7[1]), .B0(d7[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[2]), .B1(d7[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16223), .COUT(n16224), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[0]), .B1(d7[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16223), .S1(d8_71__N_1603[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1592_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_38 (.A0(d_d_tmp[71]), .B0(d_tmp[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16222), .S0(n78_adj_5051));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1550_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_36 (.A0(d_d_tmp[69]), .B0(d_tmp[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[70]), .B1(d_tmp[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16221), .COUT(n16222), .S0(n84_adj_5053), 
          .S1(n81_adj_5052));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_34 (.A0(d_d_tmp[67]), .B0(d_tmp[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[68]), .B1(d_tmp[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16220), .COUT(n16221), .S0(n90_adj_5055), 
          .S1(n87_adj_5054));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_32 (.A0(d_d_tmp[65]), .B0(d_tmp[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[66]), .B1(d_tmp[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16219), .COUT(n16220), .S0(n96_adj_5057), 
          .S1(n93_adj_5056));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_30 (.A0(d_d_tmp[63]), .B0(d_tmp[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[64]), .B1(d_tmp[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16218), .COUT(n16219), .S0(n102_adj_5059), 
          .S1(n99_adj_5058));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_28 (.A0(d_d_tmp[61]), .B0(d_tmp[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[62]), .B1(d_tmp[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16217), .COUT(n16218), .S0(n108_adj_5061), 
          .S1(n105_adj_5060));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_26 (.A0(d_d_tmp[59]), .B0(d_tmp[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[60]), .B1(d_tmp[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16216), .COUT(n16217), .S0(n114_adj_5063), 
          .S1(n111_adj_5062));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_24 (.A0(d_d_tmp[57]), .B0(d_tmp[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[58]), .B1(d_tmp[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16215), .COUT(n16216), .S0(n120_adj_5065), 
          .S1(n117_adj_5064));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_22 (.A0(d_d_tmp[55]), .B0(d_tmp[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[56]), .B1(d_tmp[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16214), .COUT(n16215), .S0(n126_adj_5067), 
          .S1(n123_adj_5066));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_20 (.A0(d_d_tmp[53]), .B0(d_tmp[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[54]), .B1(d_tmp[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16213), .COUT(n16214), .S0(n132_adj_5069), 
          .S1(n129_adj_5068));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_18 (.A0(d_d_tmp[51]), .B0(d_tmp[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[52]), .B1(d_tmp[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16212), .COUT(n16213), .S0(n138_adj_5071), 
          .S1(n135_adj_5070));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_16 (.A0(d_d_tmp[49]), .B0(d_tmp[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[50]), .B1(d_tmp[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16211), .COUT(n16212), .S0(n144_adj_5073), 
          .S1(n141_adj_5072));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_14 (.A0(d_d_tmp[47]), .B0(d_tmp[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[48]), .B1(d_tmp[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16210), .COUT(n16211), .S0(n150_adj_5075), 
          .S1(n147_adj_5074));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_12 (.A0(d_d_tmp[45]), .B0(d_tmp[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[46]), .B1(d_tmp[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16209), .COUT(n16210), .S0(n156_adj_5077), 
          .S1(n153_adj_5076));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_10 (.A0(d_d_tmp[43]), .B0(d_tmp[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[44]), .B1(d_tmp[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16208), .COUT(n16209), .S0(n162_adj_5079), 
          .S1(n159_adj_5078));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_8 (.A0(d_d_tmp[41]), .B0(d_tmp[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[42]), .B1(d_tmp[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16207), .COUT(n16208), .S0(n168_adj_5081), 
          .S1(n165_adj_5080));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_6 (.A0(d_d_tmp[39]), .B0(d_tmp[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[40]), .B1(d_tmp[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16206), .COUT(n16207), .S0(n174_adj_5083), 
          .S1(n171_adj_5082));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_4 (.A0(d_d_tmp[37]), .B0(d_tmp[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[38]), .B1(d_tmp[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16205), .COUT(n16206), .S0(n180_adj_5085), 
          .S1(n177_adj_5084));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1550_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[36]), .B1(d_tmp[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16205), .S1(n183_adj_5086));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1550_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1550_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1550_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_38 (.A0(d_d7[71]), .B0(d7[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16204), .S0(n78_adj_4924));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1640_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_36 (.A0(d_d7[69]), .B0(d7[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[70]), .B1(d7[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16203), .COUT(n16204), .S0(n84_adj_4926), .S1(n81_adj_4925));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_34 (.A0(d_d7[67]), .B0(d7[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[68]), .B1(d7[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16202), .COUT(n16203), .S0(n90_adj_4928), .S1(n87_adj_4927));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_32 (.A0(d_d7[65]), .B0(d7[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[66]), .B1(d7[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16201), .COUT(n16202), .S0(n96_adj_4930), .S1(n93_adj_4929));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_30 (.A0(d_d7[63]), .B0(d7[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[64]), .B1(d7[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16200), .COUT(n16201), .S0(n102_adj_4932), .S1(n99_adj_4931));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_28 (.A0(d_d7[61]), .B0(d7[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[62]), .B1(d7[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16199), .COUT(n16200), .S0(n108_adj_4934), .S1(n105_adj_4933));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_26 (.A0(d_d7[59]), .B0(d7[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[60]), .B1(d7[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16198), .COUT(n16199), .S0(n114_adj_4936), .S1(n111_adj_4935));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_24 (.A0(d_d7[57]), .B0(d7[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[58]), .B1(d7[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16197), .COUT(n16198), .S0(n120_adj_4938), .S1(n117_adj_4937));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_22 (.A0(d_d7[55]), .B0(d7[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[56]), .B1(d7[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16196), .COUT(n16197), .S0(n126_adj_4940), .S1(n123_adj_4939));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_20 (.A0(d_d7[53]), .B0(d7[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[54]), .B1(d7[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16195), .COUT(n16196), .S0(n132_adj_4942), .S1(n129_adj_4941));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_18 (.A0(d_d7[51]), .B0(d7[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[52]), .B1(d7[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16194), .COUT(n16195), .S0(n138_adj_4944), .S1(n135_adj_4943));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_16 (.A0(d_d7[49]), .B0(d7[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[50]), .B1(d7[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16193), .COUT(n16194), .S0(n144_adj_4946), .S1(n141_adj_4945));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_14 (.A0(d_d7[47]), .B0(d7[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[48]), .B1(d7[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16192), .COUT(n16193), .S0(n150_adj_4948), .S1(n147_adj_4947));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_12 (.A0(d_d7[45]), .B0(d7[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[46]), .B1(d7[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16191), .COUT(n16192), .S0(n156_adj_4950), .S1(n153_adj_4949));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_10 (.A0(d_d7[43]), .B0(d7[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[44]), .B1(d7[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16190), .COUT(n16191), .S0(n162_adj_4952), .S1(n159_adj_4951));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_8 (.A0(d_d7[41]), .B0(d7[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[42]), .B1(d7[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16189), .COUT(n16190), .S0(n168_adj_4954), .S1(n165_adj_4953));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_6 (.A0(d_d7[39]), .B0(d7[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[40]), .B1(d7[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16188), .COUT(n16189), .S0(n174_adj_4956), .S1(n171_adj_4955));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_4 (.A0(d_d7[37]), .B0(d7[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[38]), .B1(d7[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16187), .COUT(n16188), .S0(n180_adj_4958), .S1(n177_adj_4957));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[36]), .B1(d7[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16187), .S1(n183_adj_4959));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam _add_1_1640_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1640_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_38 (.A0(d_d6[71]), .B0(d6[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16186), .S0(n78_adj_4960));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1643_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_36 (.A0(d_d6[69]), .B0(d6[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[70]), .B1(d6[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16185), .COUT(n16186), .S0(n84_adj_4962), .S1(n81_adj_4961));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_34 (.A0(d_d6[67]), .B0(d6[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[68]), .B1(d6[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16184), .COUT(n16185), .S0(n90_adj_4964), .S1(n87_adj_4963));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_32 (.A0(d_d6[65]), .B0(d6[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[66]), .B1(d6[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16183), .COUT(n16184), .S0(n96_adj_4966), .S1(n93_adj_4965));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_30 (.A0(d_d6[63]), .B0(d6[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[64]), .B1(d6[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16182), .COUT(n16183), .S0(n102_adj_4968), .S1(n99_adj_4967));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_28 (.A0(d_d6[61]), .B0(d6[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[62]), .B1(d6[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16181), .COUT(n16182), .S0(n108_adj_4970), .S1(n105_adj_4969));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_26 (.A0(d_d6[59]), .B0(d6[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[60]), .B1(d6[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16180), .COUT(n16181), .S0(n114_adj_4972), .S1(n111_adj_4971));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_24 (.A0(d_d6[57]), .B0(d6[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[58]), .B1(d6[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16179), .COUT(n16180), .S0(n120_adj_4974), .S1(n117_adj_4973));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_22 (.A0(d_d6[55]), .B0(d6[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[56]), .B1(d6[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16178), .COUT(n16179), .S0(n126_adj_4976), .S1(n123_adj_4975));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_20 (.A0(d_d6[53]), .B0(d6[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[54]), .B1(d6[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16177), .COUT(n16178), .S0(n132_adj_4978), .S1(n129_adj_4977));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_18 (.A0(d_d6[51]), .B0(d6[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[52]), .B1(d6[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16176), .COUT(n16177), .S0(n138_adj_4980), .S1(n135_adj_4979));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_16 (.A0(d_d6[49]), .B0(d6[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[50]), .B1(d6[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16175), .COUT(n16176), .S0(n144_adj_4982), .S1(n141_adj_4981));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_14 (.A0(d_d6[47]), .B0(d6[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[48]), .B1(d6[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16174), .COUT(n16175), .S0(n150_adj_4984), .S1(n147_adj_4983));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_12 (.A0(d_d6[45]), .B0(d6[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[46]), .B1(d6[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16173), .COUT(n16174), .S0(n156_adj_4986), .S1(n153_adj_4985));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_10 (.A0(d_d6[43]), .B0(d6[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[44]), .B1(d6[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16172), .COUT(n16173), .S0(n162_adj_4988), .S1(n159_adj_4987));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_8 (.A0(d_d6[41]), .B0(d6[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[42]), .B1(d6[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16171), .COUT(n16172), .S0(n168_adj_4990), .S1(n165_adj_4989));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_6 (.A0(d_d6[39]), .B0(d6[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[40]), .B1(d6[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16170), .COUT(n16171), .S0(n174_adj_4992), .S1(n171_adj_4991));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_4 (.A0(d_d6[37]), .B0(d6[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[38]), .B1(d6[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16169), .COUT(n16170), .S0(n180_adj_4994), .S1(n177_adj_4993));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[36]), .B1(d6[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16169), .S1(n183_adj_4995));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1643_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1643_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_61 (.A0(phase_inc_carrGen[63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16168), .S0(n124));
    defparam _add_1_1412_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_1412_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_59 (.A0(phase_inc_carrGen[61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16167), .COUT(n16168), .S0(n130), 
          .S1(n127));
    defparam _add_1_1412_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_57 (.A0(phase_inc_carrGen[59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16166), .COUT(n16167), .S0(n136), 
          .S1(n133));
    defparam _add_1_1412_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_55 (.A0(phase_inc_carrGen[57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16165), .COUT(n16166), .S0(n142), 
          .S1(n139));
    defparam _add_1_1412_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_53 (.A0(phase_inc_carrGen[55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16164), .COUT(n16165), .S0(n148), 
          .S1(n145));
    defparam _add_1_1412_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_51 (.A0(phase_inc_carrGen[53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16163), .COUT(n16164), .S0(n154), 
          .S1(n151));
    defparam _add_1_1412_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_49 (.A0(phase_inc_carrGen[51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16162), .COUT(n16163), .S0(n160), 
          .S1(n157));
    defparam _add_1_1412_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_47 (.A0(phase_inc_carrGen[49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16161), .COUT(n16162), .S0(n166), 
          .S1(n163));
    defparam _add_1_1412_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_45 (.A0(phase_inc_carrGen[47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16160), .COUT(n16161), .S0(n172), 
          .S1(n169));
    defparam _add_1_1412_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_43 (.A0(phase_inc_carrGen[45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16159), .COUT(n16160), .S0(n178), 
          .S1(n175));
    defparam _add_1_1412_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_41 (.A0(phase_inc_carrGen[43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16158), .COUT(n16159), .S0(n184), 
          .S1(n181));
    defparam _add_1_1412_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_39 (.A0(phase_inc_carrGen[41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16157), .COUT(n16158), .S0(n190), 
          .S1(n187));
    defparam _add_1_1412_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_37 (.A0(phase_inc_carrGen[39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16156), .COUT(n16157), .S0(n196), 
          .S1(n193));
    defparam _add_1_1412_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_35 (.A0(phase_inc_carrGen[37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16155), .COUT(n16156), .S0(n202), 
          .S1(n199));
    defparam _add_1_1412_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_33 (.A0(phase_inc_carrGen[35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16154), .COUT(n16155), .S0(n208), 
          .S1(n205));
    defparam _add_1_1412_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_31 (.A0(phase_inc_carrGen[33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16153), .COUT(n16154), .S0(n214), 
          .S1(n211));
    defparam _add_1_1412_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_29 (.A0(phase_inc_carrGen[31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16152), .COUT(n16153), .S0(n220), 
          .S1(n217));
    defparam _add_1_1412_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_27 (.A0(phase_inc_carrGen[29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16151), .COUT(n16152), .S0(n226), 
          .S1(n223));
    defparam _add_1_1412_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_25 (.A0(phase_inc_carrGen[27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16150), .COUT(n16151), .S0(n232), 
          .S1(n229));
    defparam _add_1_1412_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_23 (.A0(phase_inc_carrGen[25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16149), .COUT(n16150), .S0(n238), 
          .S1(n235));
    defparam _add_1_1412_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_21 (.A0(phase_inc_carrGen[23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16148), .COUT(n16149), .S0(n244), 
          .S1(n241));
    defparam _add_1_1412_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_19 (.A0(phase_inc_carrGen[21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16147), .COUT(n16148), .S0(n250), 
          .S1(n247));
    defparam _add_1_1412_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_17 (.A0(phase_inc_carrGen[19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16146), .COUT(n16147), .S0(n256), 
          .S1(n253));
    defparam _add_1_1412_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_15 (.A0(phase_inc_carrGen[17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16145), .COUT(n16146), .S0(n262), 
          .S1(n259));
    defparam _add_1_1412_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_13 (.A0(phase_inc_carrGen[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16144), .COUT(n16145), .S0(n268), 
          .S1(n265));
    defparam _add_1_1412_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_11 (.A0(phase_inc_carrGen[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16143), .COUT(n16144), .S0(n274), 
          .S1(n271));
    defparam _add_1_1412_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_9 (.A0(phase_inc_carrGen[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16142), .COUT(n16143), .S0(n280), 
          .S1(n277));
    defparam _add_1_1412_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_7 (.A0(phase_inc_carrGen[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16141), .COUT(n16142), .S0(n286), 
          .S1(n283));
    defparam _add_1_1412_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_5 (.A0(phase_inc_carrGen[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16140), .COUT(n16141), .S0(n292), 
          .S1(n289));
    defparam _add_1_1412_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_3 (.A0(phase_inc_carrGen[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16139), .COUT(n16140), .S0(n298), 
          .S1(n295));
    defparam _add_1_1412_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16139), .S1(n301));
    defparam _add_1_1412_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1412_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_12 (.A0(counter[9]), .B0(DataInReg[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16138), .S1(cout_adj_4997));
    defparam _add_1_1649_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_12.INIT1 = 16'h0000;
    defparam _add_1_1649_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_10 (.A0(counter[7]), .B0(DataInReg[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(DataInReg[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16137), .COUT(n16138));
    defparam _add_1_1649_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_8 (.A0(counter[5]), .B0(DataInReg[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(DataInReg[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16136), .COUT(n16137));
    defparam _add_1_1649_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_6 (.A0(counter[3]), .B0(DataInReg[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(DataInReg[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16135), .COUT(n16136));
    defparam _add_1_1649_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_4 (.A0(counter[1]), .B0(DataInReg[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(DataInReg[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16134), .COUT(n16135));
    defparam _add_1_1649_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[0]), .B1(DataInReg[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16134));
    defparam _add_1_1649_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1649_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_13 (.A0(LOSine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16133), .S0(MixerOutSin_11__N_236[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1454_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_11 (.A0(LOSine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16132), .COUT(n16133), .S0(MixerOutSin_11__N_236[9]), 
          .S1(MixerOutSin_11__N_236[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_9 (.A0(LOSine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16131), .COUT(n16132), .S0(MixerOutSin_11__N_236[7]), 
          .S1(MixerOutSin_11__N_236[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_7 (.A0(LOSine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16130), .COUT(n16131), .S0(MixerOutSin_11__N_236[5]), 
          .S1(MixerOutSin_11__N_236[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_5 (.A0(LOSine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16129), .COUT(n16130), .S0(MixerOutSin_11__N_236[3]), 
          .S1(MixerOutSin_11__N_236[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_3 (.A0(LOSine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16128), .COUT(n16129), .S0(MixerOutSin_11__N_236[1]), 
          .S1(MixerOutSin_11__N_236[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16128), .S1(MixerOutSin_11__N_236[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1454_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1454_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_38 (.A0(d_d_tmp_adj_5672[35]), .B0(d_tmp_adj_5671[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16127), .S0(d6_71__N_1459_adj_5705[35]), 
          .S1(cout_adj_5489));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1613_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_36 (.A0(d_d_tmp_adj_5672[33]), .B0(d_tmp_adj_5671[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[34]), .B1(d_tmp_adj_5671[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16126), .COUT(n16127), .S0(d6_71__N_1459_adj_5705[33]), 
          .S1(d6_71__N_1459_adj_5705[34]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_34 (.A0(d_d_tmp_adj_5672[31]), .B0(d_tmp_adj_5671[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[32]), .B1(d_tmp_adj_5671[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16125), .COUT(n16126), .S0(d6_71__N_1459_adj_5705[31]), 
          .S1(d6_71__N_1459_adj_5705[32]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_32 (.A0(d_d_tmp_adj_5672[29]), .B0(d_tmp_adj_5671[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[30]), .B1(d_tmp_adj_5671[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16124), .COUT(n16125), .S0(d6_71__N_1459_adj_5705[29]), 
          .S1(d6_71__N_1459_adj_5705[30]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_30 (.A0(d_d_tmp_adj_5672[27]), .B0(d_tmp_adj_5671[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[28]), .B1(d_tmp_adj_5671[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16123), .COUT(n16124), .S0(d6_71__N_1459_adj_5705[27]), 
          .S1(d6_71__N_1459_adj_5705[28]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_28 (.A0(d_d_tmp_adj_5672[25]), .B0(d_tmp_adj_5671[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[26]), .B1(d_tmp_adj_5671[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16122), .COUT(n16123), .S0(d6_71__N_1459_adj_5705[25]), 
          .S1(d6_71__N_1459_adj_5705[26]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_26 (.A0(d_d_tmp_adj_5672[23]), .B0(d_tmp_adj_5671[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[24]), .B1(d_tmp_adj_5671[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16121), .COUT(n16122), .S0(d6_71__N_1459_adj_5705[23]), 
          .S1(d6_71__N_1459_adj_5705[24]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_24 (.A0(d_d_tmp_adj_5672[21]), .B0(d_tmp_adj_5671[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[22]), .B1(d_tmp_adj_5671[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16120), .COUT(n16121), .S0(d6_71__N_1459_adj_5705[21]), 
          .S1(d6_71__N_1459_adj_5705[22]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_22 (.A0(d_d_tmp_adj_5672[19]), .B0(d_tmp_adj_5671[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[20]), .B1(d_tmp_adj_5671[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16119), .COUT(n16120), .S0(d6_71__N_1459_adj_5705[19]), 
          .S1(d6_71__N_1459_adj_5705[20]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_20 (.A0(d_d_tmp_adj_5672[17]), .B0(d_tmp_adj_5671[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[18]), .B1(d_tmp_adj_5671[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16118), .COUT(n16119), .S0(d6_71__N_1459_adj_5705[17]), 
          .S1(d6_71__N_1459_adj_5705[18]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_18 (.A0(d_d_tmp_adj_5672[15]), .B0(d_tmp_adj_5671[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[16]), .B1(d_tmp_adj_5671[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16117), .COUT(n16118), .S0(d6_71__N_1459_adj_5705[15]), 
          .S1(d6_71__N_1459_adj_5705[16]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_16 (.A0(d_d_tmp_adj_5672[13]), .B0(d_tmp_adj_5671[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[14]), .B1(d_tmp_adj_5671[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16116), .COUT(n16117), .S0(d6_71__N_1459_adj_5705[13]), 
          .S1(d6_71__N_1459_adj_5705[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_14 (.A0(d_d_tmp_adj_5672[11]), .B0(d_tmp_adj_5671[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[12]), .B1(d_tmp_adj_5671[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16115), .COUT(n16116), .S0(d6_71__N_1459_adj_5705[11]), 
          .S1(d6_71__N_1459_adj_5705[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_12 (.A0(d_d_tmp_adj_5672[9]), .B0(d_tmp_adj_5671[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[10]), .B1(d_tmp_adj_5671[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16114), .COUT(n16115), .S0(d6_71__N_1459_adj_5705[9]), 
          .S1(d6_71__N_1459_adj_5705[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_10 (.A0(d_d_tmp_adj_5672[7]), .B0(d_tmp_adj_5671[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[8]), .B1(d_tmp_adj_5671[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16113), .COUT(n16114), .S0(d6_71__N_1459_adj_5705[7]), 
          .S1(d6_71__N_1459_adj_5705[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_8 (.A0(d_d_tmp_adj_5672[5]), .B0(d_tmp_adj_5671[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[6]), .B1(d_tmp_adj_5671[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16112), .COUT(n16113), .S0(d6_71__N_1459_adj_5705[5]), 
          .S1(d6_71__N_1459_adj_5705[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_6 (.A0(d_d_tmp_adj_5672[3]), .B0(d_tmp_adj_5671[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[4]), .B1(d_tmp_adj_5671[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16111), .COUT(n16112), .S0(d6_71__N_1459_adj_5705[3]), 
          .S1(d6_71__N_1459_adj_5705[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_4 (.A0(d_d_tmp_adj_5672[1]), .B0(d_tmp_adj_5671[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5672[2]), .B1(d_tmp_adj_5671[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16110), .COUT(n16111), .S0(d6_71__N_1459_adj_5705[1]), 
          .S1(d6_71__N_1459_adj_5705[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5672[0]), .B1(d_tmp_adj_5671[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16110), .S1(d6_71__N_1459_adj_5705[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1613_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_38 (.A0(d_d9[35]), .B0(d9[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16109), .S1(cout_adj_5612));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1619_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_36 (.A0(d_d9[33]), .B0(d9[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[34]), .B1(d9[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16108), .COUT(n16109));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_34 (.A0(d_d9[31]), .B0(d9[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[32]), .B1(d9[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16107), .COUT(n16108));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_32 (.A0(d_d9[29]), .B0(d9[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[30]), .B1(d9[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16106), .COUT(n16107));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_30 (.A0(d_d9[27]), .B0(d9[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[28]), .B1(d9[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16105), .COUT(n16106));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_28 (.A0(d_d9[25]), .B0(d9[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[26]), .B1(d9[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16104), .COUT(n16105));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_26 (.A0(d_d9[23]), .B0(d9[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[24]), .B1(d9[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16103), .COUT(n16104));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_24 (.A0(d_d9[21]), .B0(d9[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[22]), .B1(d9[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16102), .COUT(n16103));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_22 (.A0(d_d9[19]), .B0(d9[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[20]), .B1(d9[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16101), .COUT(n16102));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_53 (.A0(phase_inc_carrGen[52]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16657), .COUT(n16658), .S0(n163_adj_5401), 
          .S1(n160_adj_5400));
    defparam _add_1_1457_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_51 (.A0(phase_inc_carrGen[50]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16656), .COUT(n16657), .S0(n169_adj_5403), 
          .S1(n166_adj_5402));
    defparam _add_1_1457_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_49 (.A0(phase_inc_carrGen[48]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16655), .COUT(n16656), .S0(n175_adj_5405), 
          .S1(n172_adj_5404));
    defparam _add_1_1457_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_47 (.A0(phase_inc_carrGen[46]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16654), .COUT(n16655), .S0(n181_adj_5407), 
          .S1(n178_adj_5406));
    defparam _add_1_1457_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_45 (.A0(phase_inc_carrGen[44]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16653), .COUT(n16654), .S0(n187_adj_5409), 
          .S1(n184_adj_5408));
    defparam _add_1_1457_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_45.INJECT1_1 = "NO";
    LUT4 i5657_2_lut (.A(d4_adj_5676[0]), .B(d3_adj_5675[0]), .Z(d4_71__N_634_adj_5692[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5657_2_lut.init = 16'h6666;
    CCU2C _add_1_1457_add_4_43 (.A0(phase_inc_carrGen[42]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16652), .COUT(n16653), .S0(n193_adj_5411), 
          .S1(n190_adj_5410));
    defparam _add_1_1457_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_41 (.A0(phase_inc_carrGen[40]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16651), .COUT(n16652), .S0(n199_adj_5413), 
          .S1(n196_adj_5412));
    defparam _add_1_1457_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_39 (.A0(phase_inc_carrGen[38]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16650), .COUT(n16651), .S0(n205_adj_5415), 
          .S1(n202_adj_5414));
    defparam _add_1_1457_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_37 (.A0(phase_inc_carrGen[36]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16649), .COUT(n16650), .S0(n211_adj_5417), 
          .S1(n208_adj_5416));
    defparam _add_1_1457_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_37.INJECT1_1 = "NO";
    LUT4 i2492_4_lut (.A(n130_adj_5390), .B(n124), .C(led_c_3), .D(n18141), 
         .Z(n12223)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2492_4_lut.init = 16'hcac0;
    CCU2C _add_1_1457_add_4_35 (.A0(phase_inc_carrGen[34]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16648), .COUT(n16649), .S0(n217_adj_5419), 
          .S1(n214_adj_5418));
    defparam _add_1_1457_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_33 (.A0(phase_inc_carrGen[32]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16647), .COUT(n16648), .S0(n223_adj_5421), 
          .S1(n220_adj_5420));
    defparam _add_1_1457_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_31 (.A0(phase_inc_carrGen[30]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16646), .COUT(n16647), .S0(n229_adj_5423), 
          .S1(n226_adj_5422));
    defparam _add_1_1457_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_29 (.A0(phase_inc_carrGen[28]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16645), .COUT(n16646), .S0(n235_adj_5425), 
          .S1(n232_adj_5424));
    defparam _add_1_1457_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_27 (.A0(phase_inc_carrGen[26]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16644), .COUT(n16645), .S0(n241_adj_5427), 
          .S1(n238_adj_5426));
    defparam _add_1_1457_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_25 (.A0(phase_inc_carrGen[24]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16643), .COUT(n16644), .S0(n247_adj_5429), 
          .S1(n244_adj_5428));
    defparam _add_1_1457_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_23 (.A0(phase_inc_carrGen[22]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16642), .COUT(n16643), .S0(n253_adj_5431), 
          .S1(n250_adj_5430));
    defparam _add_1_1457_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_21 (.A0(phase_inc_carrGen[20]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16641), .COUT(n16642), .S0(n259_adj_5433), 
          .S1(n256_adj_5432));
    defparam _add_1_1457_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_19 (.A0(phase_inc_carrGen[18]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16640), .COUT(n16641), .S0(n265_adj_5435), 
          .S1(n262_adj_5434));
    defparam _add_1_1457_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_17 (.A0(phase_inc_carrGen[16]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16639), .COUT(n16640), .S0(n271_adj_5437), 
          .S1(n268_adj_5436));
    defparam _add_1_1457_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_15 (.A0(phase_inc_carrGen[14]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16638), .COUT(n16639), .S0(n277_adj_5439), 
          .S1(n274_adj_5438));
    defparam _add_1_1457_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_13 (.A0(phase_inc_carrGen[12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16637), .COUT(n16638), .S0(n283_adj_5441), 
          .S1(n280_adj_5440));
    defparam _add_1_1457_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_1457_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_11 (.A0(phase_inc_carrGen[10]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16636), .COUT(n16637), .S0(n289_adj_5443), 
          .S1(n286_adj_5442));
    defparam _add_1_1457_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_9 (.A0(phase_inc_carrGen[8]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16635), .COUT(n16636), .S0(n295_adj_5445), 
          .S1(n292_adj_5444));
    defparam _add_1_1457_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_7 (.A0(phase_inc_carrGen[6]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16634), .COUT(n16635), .S0(n301_adj_5447), 
          .S1(n298_adj_5446));
    defparam _add_1_1457_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_5 (.A0(phase_inc_carrGen[4]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16633), .COUT(n16634), .S0(n307), 
          .S1(n304));
    defparam _add_1_1457_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_3 (.A0(phase_inc_carrGen[2]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[3]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16632), .COUT(n16633), .S0(n313), 
          .S1(n310));
    defparam _add_1_1457_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1457_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1457_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16632), .S1(n316));
    defparam _add_1_1457_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1457_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1457_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_1.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_64 (.A0(phase_inc_carrGen1[62]), .B0(phase_accum[62]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[63]), .B1(phase_accum[63]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16630), .S0(n135_adj_4786), 
          .S1(n132_adj_4787));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_64.INIT0 = 16'h666a;
    defparam phase_accum_add_4_64.INIT1 = 16'h666a;
    defparam phase_accum_add_4_64.INJECT1_0 = "NO";
    defparam phase_accum_add_4_64.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_62 (.A0(phase_inc_carrGen1[60]), .B0(phase_accum[60]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[61]), .B1(phase_accum[61]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16629), .COUT(n16630), .S0(n141_adj_4784), 
          .S1(n138_adj_4785));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_62.INIT0 = 16'h666a;
    defparam phase_accum_add_4_62.INIT1 = 16'h666a;
    defparam phase_accum_add_4_62.INJECT1_0 = "NO";
    defparam phase_accum_add_4_62.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_60 (.A0(phase_inc_carrGen1[58]), .B0(phase_accum[58]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[59]), .B1(phase_accum[59]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16628), .COUT(n16629), .S0(n147_adj_4754), 
          .S1(n144_adj_4769));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_60.INIT0 = 16'h666a;
    defparam phase_accum_add_4_60.INIT1 = 16'h666a;
    defparam phase_accum_add_4_60.INJECT1_0 = "NO";
    defparam phase_accum_add_4_60.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_58 (.A0(phase_inc_carrGen1[56]), .B0(phase_accum[56]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[57]), .B1(phase_accum[57]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16627), .COUT(n16628), .S0(n153_adj_4752), 
          .S1(n150_adj_4753));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_58.INIT0 = 16'h666a;
    defparam phase_accum_add_4_58.INIT1 = 16'h666a;
    defparam phase_accum_add_4_58.INJECT1_0 = "NO";
    defparam phase_accum_add_4_58.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_56 (.A0(phase_inc_carrGen1[54]), .B0(phase_accum_adj_5665[54]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[55]), .B1(phase_accum_adj_5665[55]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16626), .COUT(n16627), .S0(n159_adj_4750), 
          .S1(n156_adj_4751));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_56.INIT0 = 16'h666a;
    defparam phase_accum_add_4_56.INIT1 = 16'h666a;
    defparam phase_accum_add_4_56.INJECT1_0 = "NO";
    defparam phase_accum_add_4_56.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_54 (.A0(phase_inc_carrGen1[52]), .B0(phase_accum_adj_5665[52]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[53]), .B1(phase_accum_adj_5665[53]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16625), .COUT(n16626), .S0(n165_adj_4748), 
          .S1(n162_adj_4749));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_54.INIT0 = 16'h666a;
    defparam phase_accum_add_4_54.INIT1 = 16'h666a;
    defparam phase_accum_add_4_54.INJECT1_0 = "NO";
    defparam phase_accum_add_4_54.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_52 (.A0(phase_inc_carrGen1[50]), .B0(phase_accum_adj_5665[50]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[51]), .B1(phase_accum_adj_5665[51]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16624), .COUT(n16625), .S0(n171_adj_4738), 
          .S1(n168_adj_4743));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_52.INIT0 = 16'h666a;
    defparam phase_accum_add_4_52.INIT1 = 16'h666a;
    defparam phase_accum_add_4_52.INJECT1_0 = "NO";
    defparam phase_accum_add_4_52.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_50 (.A0(phase_inc_carrGen1[48]), .B0(phase_accum_adj_5665[48]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[49]), .B1(phase_accum_adj_5665[49]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16623), .COUT(n16624), .S0(n177_adj_4735), 
          .S1(n174_adj_4737));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_50.INIT0 = 16'h666a;
    defparam phase_accum_add_4_50.INIT1 = 16'h666a;
    defparam phase_accum_add_4_50.INJECT1_0 = "NO";
    defparam phase_accum_add_4_50.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_48 (.A0(phase_inc_carrGen1[46]), .B0(phase_accum_adj_5665[46]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[47]), .B1(phase_accum_adj_5665[47]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16622), .COUT(n16623), .S0(n183_adj_4733), 
          .S1(n180_adj_4734));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_48.INIT0 = 16'h666a;
    defparam phase_accum_add_4_48.INIT1 = 16'h666a;
    defparam phase_accum_add_4_48.INJECT1_0 = "NO";
    defparam phase_accum_add_4_48.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_46 (.A0(phase_inc_carrGen1[44]), .B0(phase_accum_adj_5665[44]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[45]), .B1(phase_accum_adj_5665[45]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16621), .COUT(n16622), .S0(n189), 
          .S1(n186));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_46.INIT0 = 16'h666a;
    defparam phase_accum_add_4_46.INIT1 = 16'h666a;
    defparam phase_accum_add_4_46.INJECT1_0 = "NO";
    defparam phase_accum_add_4_46.INJECT1_1 = "NO";
    LUT4 i3173_2_lut_rep_161 (.A(led_c_4), .B(n2845), .Z(n18131)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3173_2_lut_rep_161.init = 16'h8888;
    CCU2C phase_accum_add_4_44 (.A0(phase_inc_carrGen1[42]), .B0(phase_accum_adj_5665[42]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[43]), .B1(phase_accum_adj_5665[43]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16620), .COUT(n16621), .S0(n195), 
          .S1(n192));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_44.INIT0 = 16'h666a;
    defparam phase_accum_add_4_44.INIT1 = 16'h666a;
    defparam phase_accum_add_4_44.INJECT1_0 = "NO";
    defparam phase_accum_add_4_44.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_42 (.A0(phase_inc_carrGen1[40]), .B0(phase_accum_adj_5665[40]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[41]), .B1(phase_accum_adj_5665[41]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16619), .COUT(n16620), .S0(n201), 
          .S1(n198));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_42.INIT0 = 16'h666a;
    defparam phase_accum_add_4_42.INIT1 = 16'h666a;
    defparam phase_accum_add_4_42.INJECT1_0 = "NO";
    defparam phase_accum_add_4_42.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_40 (.A0(phase_inc_carrGen1[38]), .B0(phase_accum_adj_5665[38]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[39]), .B1(phase_accum_adj_5665[39]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16618), .COUT(n16619), .S0(n207), 
          .S1(n204));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_40.INIT0 = 16'h666a;
    defparam phase_accum_add_4_40.INIT1 = 16'h666a;
    defparam phase_accum_add_4_40.INJECT1_0 = "NO";
    defparam phase_accum_add_4_40.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_38 (.A0(phase_inc_carrGen1[36]), .B0(phase_accum_adj_5665[36]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[37]), .B1(phase_accum_adj_5665[37]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16617), .COUT(n16618), .S0(n213), 
          .S1(n210));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_38.INIT0 = 16'h666a;
    defparam phase_accum_add_4_38.INIT1 = 16'h666a;
    defparam phase_accum_add_4_38.INJECT1_0 = "NO";
    defparam phase_accum_add_4_38.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_36 (.A0(phase_inc_carrGen1[34]), .B0(phase_accum_adj_5665[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[35]), .B1(phase_accum_adj_5665[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16616), .COUT(n16617), .S0(n219), 
          .S1(n216));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_36.INIT0 = 16'h666a;
    defparam phase_accum_add_4_36.INIT1 = 16'h666a;
    defparam phase_accum_add_4_36.INJECT1_0 = "NO";
    defparam phase_accum_add_4_36.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_34 (.A0(phase_inc_carrGen1[32]), .B0(phase_accum_adj_5665[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[33]), .B1(phase_accum_adj_5665[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16615), .COUT(n16616), .S0(n225), 
          .S1(n222));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_34.INIT0 = 16'h666a;
    defparam phase_accum_add_4_34.INIT1 = 16'h666a;
    defparam phase_accum_add_4_34.INJECT1_0 = "NO";
    defparam phase_accum_add_4_34.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_32 (.A0(phase_inc_carrGen1[30]), .B0(phase_accum_adj_5665[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[31]), .B1(phase_accum_adj_5665[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16614), .COUT(n16615), .S0(n231), 
          .S1(n228));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_32.INIT0 = 16'h666a;
    defparam phase_accum_add_4_32.INIT1 = 16'h666a;
    defparam phase_accum_add_4_32.INJECT1_0 = "NO";
    defparam phase_accum_add_4_32.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_30 (.A0(phase_inc_carrGen1[28]), .B0(phase_accum_adj_5665[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[29]), .B1(phase_accum_adj_5665[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16613), .COUT(n16614), .S0(n237), 
          .S1(n234));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_30.INIT0 = 16'h666a;
    defparam phase_accum_add_4_30.INIT1 = 16'h666a;
    defparam phase_accum_add_4_30.INJECT1_0 = "NO";
    defparam phase_accum_add_4_30.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_28 (.A0(phase_inc_carrGen1[26]), .B0(phase_accum_adj_5665[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[27]), .B1(phase_accum_adj_5665[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16612), .COUT(n16613), .S0(n243), 
          .S1(n240));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_28.INIT0 = 16'h666a;
    defparam phase_accum_add_4_28.INIT1 = 16'h666a;
    defparam phase_accum_add_4_28.INJECT1_0 = "NO";
    defparam phase_accum_add_4_28.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_26 (.A0(phase_inc_carrGen1[24]), .B0(phase_accum_adj_5665[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[25]), .B1(phase_accum_adj_5665[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16611), .COUT(n16612), .S0(n249), 
          .S1(n246));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_26.INIT0 = 16'h666a;
    defparam phase_accum_add_4_26.INIT1 = 16'h666a;
    defparam phase_accum_add_4_26.INJECT1_0 = "NO";
    defparam phase_accum_add_4_26.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_24 (.A0(phase_inc_carrGen1[22]), .B0(phase_accum_adj_5665[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[23]), .B1(phase_accum_adj_5665[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16610), .COUT(n16611), .S0(n255), 
          .S1(n252));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_24.INIT0 = 16'h666a;
    defparam phase_accum_add_4_24.INIT1 = 16'h666a;
    defparam phase_accum_add_4_24.INJECT1_0 = "NO";
    defparam phase_accum_add_4_24.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_22 (.A0(phase_inc_carrGen1[20]), .B0(phase_accum_adj_5665[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[21]), .B1(phase_accum_adj_5665[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16609), .COUT(n16610), .S0(n261), 
          .S1(n258));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_22.INIT0 = 16'h666a;
    defparam phase_accum_add_4_22.INIT1 = 16'h666a;
    defparam phase_accum_add_4_22.INJECT1_0 = "NO";
    defparam phase_accum_add_4_22.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_20 (.A0(phase_inc_carrGen1[18]), .B0(phase_accum_adj_5665[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[19]), .B1(phase_accum_adj_5665[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16608), .COUT(n16609), .S0(n267), 
          .S1(n264));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_20.INIT0 = 16'h666a;
    defparam phase_accum_add_4_20.INIT1 = 16'h666a;
    defparam phase_accum_add_4_20.INJECT1_0 = "NO";
    defparam phase_accum_add_4_20.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_18 (.A0(phase_inc_carrGen1[16]), .B0(phase_accum_adj_5665[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[17]), .B1(phase_accum_adj_5665[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16607), .COUT(n16608), .S0(n273), 
          .S1(n270));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_18.INIT0 = 16'h666a;
    defparam phase_accum_add_4_18.INIT1 = 16'h666a;
    defparam phase_accum_add_4_18.INJECT1_0 = "NO";
    defparam phase_accum_add_4_18.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_16 (.A0(phase_inc_carrGen1[14]), .B0(phase_accum_adj_5665[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[15]), .B1(phase_accum_adj_5665[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16606), .COUT(n16607), .S0(n279), 
          .S1(n276));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_16.INIT0 = 16'h666a;
    defparam phase_accum_add_4_16.INIT1 = 16'h666a;
    defparam phase_accum_add_4_16.INJECT1_0 = "NO";
    defparam phase_accum_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_14 (.A0(phase_inc_carrGen1[12]), .B0(phase_accum_adj_5665[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[13]), .B1(phase_accum_adj_5665[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16605), .COUT(n16606), .S0(n285), 
          .S1(n282));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_14.INIT0 = 16'h666a;
    defparam phase_accum_add_4_14.INIT1 = 16'h666a;
    defparam phase_accum_add_4_14.INJECT1_0 = "NO";
    defparam phase_accum_add_4_14.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_12 (.A0(phase_inc_carrGen1[10]), .B0(phase_accum_adj_5665[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[11]), .B1(phase_accum_adj_5665[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16604), .COUT(n16605), .S0(n291), 
          .S1(n288));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_12.INIT0 = 16'h666a;
    defparam phase_accum_add_4_12.INIT1 = 16'h666a;
    defparam phase_accum_add_4_12.INJECT1_0 = "NO";
    defparam phase_accum_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_20 (.A0(d_d9[17]), .B0(d9[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[18]), .B1(d9[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16100), .COUT(n16101));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_18 (.A0(d_d9[15]), .B0(d9[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[16]), .B1(d9[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16099), .COUT(n16100));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_16 (.A0(d_d9[13]), .B0(d9[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[14]), .B1(d9[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16098), .COUT(n16099));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_14 (.A0(d_d9[11]), .B0(d9[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[12]), .B1(d9[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16097), .COUT(n16098));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_12 (.A0(d_d9[9]), .B0(d9[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[10]), .B1(d9[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16096), .COUT(n16097));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_10 (.A0(d_d9[7]), .B0(d9[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[8]), .B1(d9[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16095), .COUT(n16096));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_8 (.A0(d_d9[5]), .B0(d9[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[6]), .B1(d9[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16094), .COUT(n16095));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_6 (.A0(d_d9[3]), .B0(d9[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[4]), .B1(d9[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16093), .COUT(n16094));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_4 (.A0(d_d9[1]), .B0(d9[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[2]), .B1(d9[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16092), .COUT(n16093));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[0]), .B1(d9[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16092));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1619_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_38 (.A0(d1_adj_5673[71]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16091), .S0(n78_adj_5576));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1568_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_36 (.A0(d1_adj_5673[69]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[70]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16090), .COUT(n16091), .S0(n84_adj_5578), 
          .S1(n81_adj_5577));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_34 (.A0(d1_adj_5673[67]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[68]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16089), .COUT(n16090), .S0(n90_adj_5580), 
          .S1(n87_adj_5579));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_32 (.A0(d1_adj_5673[65]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[66]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16088), .COUT(n16089), .S0(n96_adj_5582), 
          .S1(n93_adj_5581));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_30 (.A0(d1_adj_5673[63]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[64]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16087), .COUT(n16088), .S0(n102_adj_5584), 
          .S1(n99_adj_5583));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_28 (.A0(d1_adj_5673[61]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[62]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16086), .COUT(n16087), .S0(n108_adj_5586), 
          .S1(n105_adj_5585));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_26 (.A0(d1_adj_5673[59]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[60]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16085), .COUT(n16086), .S0(n114_adj_5588), 
          .S1(n111_adj_5587));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_24 (.A0(d1_adj_5673[57]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[58]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16084), .COUT(n16085), .S0(n120_adj_5590), 
          .S1(n117_adj_5589));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_22 (.A0(d1_adj_5673[55]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[56]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16083), .COUT(n16084), .S0(n126_adj_5592), 
          .S1(n123_adj_5591));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_20 (.A0(d1_adj_5673[53]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5673[54]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16082), .COUT(n16083), .S0(n132_adj_5594), 
          .S1(n129_adj_5593));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1568_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_20.INJECT1_1 = "NO";
    LUT4 i2250_3_lut_4_lut (.A(n18138), .B(n18267), .C(led_c_3), .D(n298), 
         .Z(n11965)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2250_3_lut_4_lut.init = 16'hf808;
    LUT4 n18075_bdd_4_lut (.A(n18075), .B(n18074), .C(led_c_0), .D(n18139), 
         .Z(n18127)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n18075_bdd_4_lut.init = 16'hffca;
    LUT4 i2322_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(led_c_3), .D(n172), 
         .Z(n12037)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2322_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_326_i61_4_lut (.A(n12059), .B(n139_adj_5393), .C(n18135), 
         .D(n2593), .Z(n2332)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i61_4_lut.init = 16'hc0ca;
    LUT4 i2488_4_lut (.A(n136_adj_5392), .B(n130), .C(led_c_3), .D(n18141), 
         .Z(n12219)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2488_4_lut.init = 16'hcac0;
    LUT4 i2306_3_lut_4_lut (.A(n18138), .B(n18267), .C(n18268), .D(n202), 
         .Z(n12021)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2306_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_326_i59_4_lut (.A(n12055), .B(n145_adj_5395), .C(n18135), 
         .D(n2593), .Z(n2334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i59_4_lut.init = 16'hcfca;
    LUT4 i5654_2_lut (.A(d5_adj_5677[0]), .B(d4_adj_5676[0]), .Z(d5_71__N_706_adj_5693[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5654_2_lut.init = 16'h6666;
    CCU2C add_4105_11 (.A0(ISquare[31]), .B0(n18150), .C0(n18143), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n18150), .C1(n18143), .D1(VCC_net), 
          .CIN(n16785), .S0(n44), .S1(d_out_d_11__N_1874[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4105_11.INIT0 = 16'he1e1;
    defparam add_4105_11.INIT1 = 16'he1e1;
    defparam add_4105_11.INJECT1_0 = "NO";
    defparam add_4105_11.INJECT1_1 = "NO";
    LUT4 i3257_1_lut_2_lut (.A(led_c_4), .B(n2845), .Z(n3685)) /* synthesis lut_function=(!(A (B))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3257_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_326_i60_4_lut (.A(n12057), .B(n142_adj_5394), .C(n18135), 
         .D(n2593), .Z(n2333)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i60_4_lut.init = 16'hc0ca;
    LUT4 mux_326_i57_4_lut (.A(n2536), .B(n151_adj_5397), .C(n18135), 
         .D(n2593), .Z(n2336)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i57_4_lut.init = 16'hc0ca;
    LUT4 i2486_4_lut (.A(n148_adj_5396), .B(n142), .C(led_c_3), .D(n18141), 
         .Z(n12217)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2486_4_lut.init = 16'hcac0;
    CCU2C add_4105_9 (.A0(n18143), .B0(ISquare[31]), .C0(ISquare[23]), 
          .D0(ISquare[22]), .A1(n40), .B1(n15364), .C1(n209), .D1(ISquare[31]), 
          .CIN(n16784), .COUT(n16785), .S0(n50), .S1(n47));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4105_9.INIT0 = 16'h6665;
    defparam add_4105_9.INIT1 = 16'h556a;
    defparam add_4105_9.INJECT1_0 = "NO";
    defparam add_4105_9.INJECT1_1 = "NO";
    LUT4 mux_326_i55_4_lut (.A(n12049), .B(n157_adj_5399), .C(n18135), 
         .D(n2593), .Z(n2338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i55_4_lut.init = 16'hcfca;
    LUT4 i1_3_lut_4_lut_4_lut (.A(led_c_0), .B(led_c_6), .C(n11_adj_4564), 
         .D(led_c_1), .Z(n17595)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.A(n18138), .B(led_c_2), .C(n18134), 
         .D(led_c_3), .Z(n17496)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_2_lut_3_lut_4_lut_adj_58.init = 16'h0008;
    CCU2C add_4105_7 (.A0(n49), .B0(ISquare[31]), .C0(ISquare[23]), .D0(ISquare[22]), 
          .A1(n18150), .B1(ISquare[31]), .C1(ISquare[23]), .D1(ISquare[22]), 
          .CIN(n16783), .COUT(n16784), .S0(n56), .S1(n53));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4105_7.INIT0 = 16'h999a;
    defparam add_4105_7.INIT1 = 16'haaa9;
    defparam add_4105_7.INJECT1_0 = "NO";
    defparam add_4105_7.INJECT1_1 = "NO";
    LUT4 mux_326_i56_4_lut (.A(n2403), .B(n154_adj_5398), .C(n18135), 
         .D(n12136), .Z(n2337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i56_4_lut.init = 16'hcfca;
    LUT4 i3253_2_lut (.A(n148), .B(n18268), .Z(n2403)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3253_2_lut.init = 16'h8888;
    CCU2C add_4105_5 (.A0(ISquare[22]), .B0(ISquare[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[23]), .B1(ISquare[22]), .C1(ISquare[31]), 
          .D1(n15364), .CIN(n16782), .COUT(n16783), .S0(n62), .S1(n59));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4105_5.INIT0 = 16'h9999;
    defparam add_4105_5.INIT1 = 16'heee1;
    defparam add_4105_5.INJECT1_0 = "NO";
    defparam add_4105_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_3_lut (.A(led_c_3), .B(led_c_0), .C(led_c_4), .Z(n17593)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h5454;
    LUT4 i3324_2_lut_2_lut (.A(led_c_3), .B(n145), .Z(n2536)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i3324_2_lut_2_lut.init = 16'hdddd;
    CCU2C add_4105_3 (.A0(ISquare[31]), .B0(n18150), .C0(ISquare[20]), 
          .D0(VCC_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16781), .COUT(n16782), .S1(n65_adj_5486));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4105_3.INIT0 = 16'he1e1;
    defparam add_4105_3.INIT1 = 16'h555f;
    defparam add_4105_3.INJECT1_0 = "NO";
    defparam add_4105_3.INJECT1_1 = "NO";
    CCU2C add_4105_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[22]), .B1(ISquare[23]), .C1(n209), .D1(ISquare[31]), 
          .COUT(n16781));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4105_1.INIT0 = 16'h0000;
    defparam add_4105_1.INIT1 = 16'h001f;
    defparam add_4105_1.INJECT1_0 = "NO";
    defparam add_4105_1.INJECT1_1 = "NO";
    LUT4 i2484_4_lut (.A(n163_adj_5401), .B(n157), .C(led_c_3), .D(n18141), 
         .Z(n12215)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2484_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_4_lut_4_lut (.A(led_c_3), .B(n18137), .C(n18144), .D(n26_adj_5659), 
         .Z(n12136)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h5400;
    LUT4 i3318_2_lut_2_lut (.A(n18268), .B(n226), .Z(n2563)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i3318_2_lut_2_lut.init = 16'hdddd;
    LUT4 led_c_0_bdd_4_lut_3_lut (.A(led_c_3), .B(n18267), .C(led_c_1), 
         .Z(n18075)) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam led_c_0_bdd_4_lut_3_lut.init = 16'h6f6f;
    LUT4 i27_3_lut_4_lut_4_lut (.A(led_c_3), .B(n193), .C(n26_adj_5659), 
         .D(n18144), .Z(n13_adj_5488)) /* synthesis lut_function=(!(A (B)+!A !(C (D)))) */ ;
    defparam i27_3_lut_4_lut_4_lut.init = 16'h7222;
    LUT4 i2316_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(n18268), .D(n184), 
         .Z(n12031)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2316_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i6134_3_lut_4_lut_4_lut (.A(led_c_3), .B(n18134), .C(n18267), 
         .D(n18138), .Z(n17322)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;
    defparam i6134_3_lut_4_lut_4_lut.init = 16'h5444;
    LUT4 i27_3_lut_4_lut_4_lut_adj_59 (.A(led_c_3), .B(n247), .C(n26_adj_5659), 
         .D(n18144), .Z(n13_adj_5485)) /* synthesis lut_function=(!(A (B)+!A !(C (D)))) */ ;
    defparam i27_3_lut_4_lut_4_lut_adj_59.init = 16'h7222;
    LUT4 i6635_4_lut (.A(led_c_2), .B(n17319), .C(led_c_3), .D(led_c_6), 
         .Z(clk_80mhz_enable_1470)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i6635_4_lut.init = 16'h0001;
    LUT4 i3251_2_lut_2_lut (.A(led_c_3), .B(n181), .Z(n2414)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i3251_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_326_i54_4_lut (.A(n12047), .B(n160_adj_5400), .C(n18135), 
         .D(n2593), .Z(n2339)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i54_4_lut.init = 16'hc0ca;
    LUT4 mux_326_i18_4_lut (.A(n2575), .B(n268_adj_5436), .C(n18135), 
         .D(n2593), .Z(n2375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i18_4_lut.init = 16'hcfca;
    LUT4 i3248_2_lut_2_lut (.A(led_c_3), .B(n268), .Z(n2443)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i3248_2_lut_2_lut.init = 16'hdddd;
    LUT4 i6595_3_lut (.A(led_c_3), .B(n18301), .C(n13099), .Z(clk_80mhz_enable_831)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;
    defparam i6595_3_lut.init = 16'hc4c4;
    LUT4 i3310_2_lut_2_lut (.A(led_c_3), .B(n295), .Z(n2586)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i3310_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2296_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(led_c_3), .D(n217), 
         .Z(n12011)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2296_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i3315_2_lut (.A(n262), .B(n18268), .Z(n2575)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3315_2_lut.init = 16'h8888;
    LUT4 mux_326_i15_4_lut (.A(n7_adj_5660), .B(n277_adj_5439), .C(n18135), 
         .D(n17322), .Z(n2378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i15_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_adj_60 (.A(n18268), .B(n271), .Z(n7_adj_5660)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_2_lut_adj_60.init = 16'h8888;
    LUT4 i2298_3_lut_4_lut (.A(n18267), .B(n18138), .C(n18268), .D(n214), 
         .Z(n12013)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2298_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_326_i16_4_lut (.A(n2443), .B(n274_adj_5438), .C(n18135), 
         .D(n12136), .Z(n2377)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i16_4_lut.init = 16'hc0ca;
    LUT4 mux_326_i13_4_lut (.A(n2446), .B(n283_adj_5441), .C(n18135), 
         .D(n12136), .Z(n2380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i13_4_lut.init = 16'hcfca;
    LUT4 i3247_2_lut (.A(n277), .B(led_c_3), .Z(n2446)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3247_2_lut.init = 16'h8888;
    LUT4 mux_326_i14_4_lut (.A(n2579), .B(n280_adj_5440), .C(n18135), 
         .D(n2593), .Z(n2379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i14_4_lut.init = 16'hcfca;
    LUT4 i3313_2_lut (.A(n274), .B(n18268), .Z(n2579)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3313_2_lut.init = 16'h8888;
    LUT4 i2280_3_lut_4_lut (.A(n18267), .B(n18138), .C(n18268), .D(n241), 
         .Z(n11995)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2280_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_326_i11_4_lut (.A(n11973), .B(n289_adj_5443), .C(n18135), 
         .D(n2593), .Z(n2382)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i11_4_lut.init = 16'hc0ca;
    LUT4 i2476_4_lut (.A(n286_adj_5442), .B(n280), .C(led_c_3), .D(n18141), 
         .Z(n12207)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2476_4_lut.init = 16'hcac0;
    LUT4 mux_326_i9_4_lut (.A(n11969), .B(n295_adj_5445), .C(n18135), 
         .D(n2593), .Z(n2384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i9_4_lut.init = 16'hcfca;
    LUT4 mux_326_i10_4_lut (.A(n11971), .B(n292_adj_5444), .C(n18135), 
         .D(n2593), .Z(n2383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i10_4_lut.init = 16'hcfca;
    LUT4 i2270_3_lut_4_lut (.A(n18267), .B(n18138), .C(led_c_3), .D(n259), 
         .Z(n11985)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2270_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_326_i7_4_lut (.A(n2586), .B(n301_adj_5447), .C(n18135), .D(n2593), 
         .Z(n2386)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i7_4_lut.init = 16'hc0ca;
    LUT4 mux_326_i8_4_lut (.A(n2451), .B(n298_adj_5446), .C(n18135), .D(n12136), 
         .Z(n2385)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i8_4_lut.init = 16'hc0ca;
    LUT4 i360_2_lut_3_lut_4_lut_4_lut (.A(led_c_3), .B(n26_adj_5659), .C(n18145), 
         .D(led_c_4), .Z(n2593)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i360_2_lut_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 mux_326_i5_4_lut (.A(n11963), .B(n307), .C(n18135), .D(n2593), 
         .Z(n2388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i5_4_lut.init = 16'hcfca;
    LUT4 mux_326_i6_4_lut (.A(n11965), .B(n304), .C(n18135), .D(n2593), 
         .Z(n2387)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i6_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1577_add_4_16 (.A0(d4_adj_5676[49]), .B0(d3_adj_5675[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[50]), .B1(d3_adj_5675[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16274), .COUT(n16275), .S0(n144_adj_4739), 
          .S1(n141_adj_4740));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_29 (.A0(d_tmp[62]), .B0(cout_adj_5496), .C0(n105_adj_5060), 
          .D0(n11_adj_4759), .A1(d_tmp[63]), .B1(cout_adj_5496), .C1(n102_adj_5059), 
          .D1(n10_adj_4760), .CIN(n16337), .COUT(n16338), .S0(d6_71__N_1459[62]), 
          .S1(d6_71__N_1459[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_29.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_10 (.A0(phase_inc_carrGen1[8]), .B0(phase_accum_adj_5665[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[9]), .B1(phase_accum_adj_5665[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16603), .COUT(n16604), .S0(n297), 
          .S1(n294));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_10.INIT0 = 16'h666a;
    defparam phase_accum_add_4_10.INIT1 = 16'h666a;
    defparam phase_accum_add_4_10.INJECT1_0 = "NO";
    defparam phase_accum_add_4_10.INJECT1_1 = "NO";
    CCU2C add_4111_13 (.A0(d_out_d_11__N_1873), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1873), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16775), .S0(n48_adj_5613), 
          .S1(d_out_d_11__N_1876[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_13.INIT0 = 16'h666a;
    defparam add_4111_13.INIT1 = 16'h666a;
    defparam add_4111_13.INJECT1_0 = "NO";
    defparam add_4111_13.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_14 (.A0(d4_adj_5676[47]), .B0(d3_adj_5675[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[48]), .B1(d3_adj_5675[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16273), .COUT(n16274), .S0(n150_adj_4562), 
          .S1(n147_adj_4563));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_14.INJECT1_1 = "NO";
    CCU2C add_4111_11 (.A0(d_out_d_11__N_1874[17]), .B0(n47), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n44), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16774), .COUT(n16775), .S0(n54_adj_5615), 
          .S1(n51_adj_5614));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_11.INIT0 = 16'h9995;
    defparam add_4111_11.INIT1 = 16'h9995;
    defparam add_4111_11.INJECT1_0 = "NO";
    defparam add_4111_11.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5685[36]), .B1(d9_adj_5684[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16495));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1637_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_2.INJECT1_1 = "NO";
    CCU2C add_4111_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1874[17]), .C0(n53), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n50), .D1(VCC_net), .CIN(n16773), .COUT(n16774), .S0(n60_adj_5617), 
          .S1(n57_adj_5616));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_9.INIT0 = 16'h6969;
    defparam add_4111_9.INIT1 = 16'h6969;
    defparam add_4111_9.INJECT1_0 = "NO";
    defparam add_4111_9.INJECT1_1 = "NO";
    CCU2C add_4111_7 (.A0(d_out_d_11__N_1874[17]), .B0(n59), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n56), .D1(VCC_net), .CIN(n16772), .COUT(n16773), .S0(n66_adj_5619), 
          .S1(n63_adj_5618));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_7.INIT0 = 16'h9995;
    defparam add_4111_7.INIT1 = 16'h6969;
    defparam add_4111_7.INJECT1_0 = "NO";
    defparam add_4111_7.INJECT1_1 = "NO";
    CCU2C add_4111_5 (.A0(n65_adj_5486), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(n18143), .C1(n62), .D1(VCC_net), 
          .CIN(n16771), .COUT(n16772), .S0(n72_adj_5621), .S1(n69_adj_5620));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_5.INIT0 = 16'haaa0;
    defparam add_4111_5.INIT1 = 16'h6969;
    defparam add_4111_5.INJECT1_0 = "NO";
    defparam add_4111_5.INJECT1_1 = "NO";
    CCU2C add_4111_3 (.A0(d_out_d_11__N_1874[17]), .B0(ISquare[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16770), .COUT(n16771), .S1(n75_adj_5622));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_3.INIT0 = 16'h666a;
    defparam add_4111_3.INIT1 = 16'h555f;
    defparam add_4111_3.INJECT1_0 = "NO";
    defparam add_4111_3.INJECT1_1 = "NO";
    CCU2C add_4111_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16770));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4111_1.INIT0 = 16'h0000;
    defparam add_4111_1.INIT1 = 16'haaaf;
    defparam add_4111_1.INJECT1_0 = "NO";
    defparam add_4111_1.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_27 (.A0(d_tmp[60]), .B0(cout_adj_5496), .C0(n111_adj_5062), 
          .D0(n13_adj_4757), .A1(d_tmp[61]), .B1(cout_adj_5496), .C1(n108_adj_5061), 
          .D1(n12_adj_4758), .CIN(n16336), .COUT(n16337), .S0(d6_71__N_1459[60]), 
          .S1(d6_71__N_1459[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_27.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_8 (.A0(phase_inc_carrGen1[6]), .B0(phase_accum_adj_5665[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[7]), .B1(phase_accum_adj_5665[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16602), .COUT(n16603), .S0(n303), 
          .S1(n300));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_8.INIT0 = 16'h666a;
    defparam phase_accum_add_4_8.INIT1 = 16'h666a;
    defparam phase_accum_add_4_8.INJECT1_0 = "NO";
    defparam phase_accum_add_4_8.INJECT1_1 = "NO";
    CCU2C add_4106_19 (.A0(d_out_d_11__N_1888[17]), .B0(n48_adj_5134), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n45_adj_5133), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16764), .S0(n45_adj_5560), 
          .S1(d_out_d_11__N_1890[17]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_19.INIT0 = 16'h9995;
    defparam add_4106_19.INIT1 = 16'h9995;
    defparam add_4106_19.INJECT1_0 = "NO";
    defparam add_4106_19.INJECT1_1 = "NO";
    CCU2C add_4106_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n54_adj_5136), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n51_adj_5135), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16763), .COUT(n16764), .S0(n51_adj_5562), 
          .S1(n48_adj_5561));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_17.INIT0 = 16'h6969;
    defparam add_4106_17.INIT1 = 16'h9995;
    defparam add_4106_17.INJECT1_0 = "NO";
    defparam add_4106_17.INJECT1_1 = "NO";
    CCU2C add_4106_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n60_adj_5138), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1888[17]), 
          .C1(n57_adj_5137), .D1(VCC_net), .CIN(n16762), .COUT(n16763), 
          .S0(n57_adj_5564), .S1(n54_adj_5563));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_15.INIT0 = 16'h6969;
    defparam add_4106_15.INIT1 = 16'h6969;
    defparam add_4106_15.INJECT1_0 = "NO";
    defparam add_4106_15.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_37 (.A0(d4_adj_5676[70]), .B0(cout_adj_5150), 
          .C0(n81_adj_4838), .D0(d5_adj_5677[70]), .A1(d4_adj_5676[71]), 
          .B1(cout_adj_5150), .C1(n78_adj_4837), .D1(d5_adj_5677[71]), 
          .CIN(n16363), .S0(d5_71__N_706_adj_5693[70]), .S1(d5_71__N_706_adj_5693[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_37.INJECT1_1 = "NO";
    CCU2C add_4106_13 (.A0(d_out_d_11__N_1888[17]), .B0(n18143), .C0(n66_adj_5140), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n63_adj_5139), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16761), .COUT(n16762), .S0(n63_adj_5566), 
          .S1(n60_adj_5565));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_13.INIT0 = 16'h6969;
    defparam add_4106_13.INIT1 = 16'h9995;
    defparam add_4106_13.INJECT1_0 = "NO";
    defparam add_4106_13.INJECT1_1 = "NO";
    CCU2C add_4106_11 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n72_adj_5142), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n69_adj_5141), .D1(VCC_net), 
          .CIN(n16760), .COUT(n16761), .S0(n69_adj_5568), .S1(n66_adj_5567));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_11.INIT0 = 16'h9696;
    defparam add_4106_11.INIT1 = 16'h9696;
    defparam add_4106_11.INJECT1_0 = "NO";
    defparam add_4106_11.INJECT1_1 = "NO";
    CCU2C add_4106_9 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n78_adj_5144), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n75_adj_5143), .D1(VCC_net), 
          .CIN(n16759), .COUT(n16760), .S0(n75_adj_5570), .S1(n72_adj_5569));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_9.INIT0 = 16'h9696;
    defparam add_4106_9.INIT1 = 16'h9696;
    defparam add_4106_9.INJECT1_0 = "NO";
    defparam add_4106_9.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_6 (.A0(phase_inc_carrGen1[4]), .B0(phase_accum_adj_5665[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[5]), .B1(phase_accum_adj_5665[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16601), .COUT(n16602), .S0(n309), 
          .S1(n306));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_6.INIT0 = 16'h666a;
    defparam phase_accum_add_4_6.INIT1 = 16'h666a;
    defparam phase_accum_add_4_6.INJECT1_0 = "NO";
    defparam phase_accum_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[36]), .B1(d3[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16535), .S1(n183_adj_5302));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1562_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_2.INJECT1_1 = "NO";
    CCU2C add_4106_7 (.A0(d_out_d_11__N_1884[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n84_adj_5146), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n81_adj_5145), .D1(VCC_net), 
          .CIN(n16758), .COUT(n16759), .S0(n81_adj_5572), .S1(n78_adj_5571));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_7.INIT0 = 16'h9696;
    defparam add_4106_7.INIT1 = 16'h9696;
    defparam add_4106_7.INJECT1_0 = "NO";
    defparam add_4106_7.INJECT1_1 = "NO";
    CCU2C add_4106_5 (.A0(n90_adj_5148), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(d_out_d_11__N_1888[17]), .C1(n87_adj_5147), 
          .D1(VCC_net), .CIN(n16757), .COUT(n16758), .S0(n87_adj_5574), 
          .S1(n84_adj_5573));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_5.INIT0 = 16'haaa0;
    defparam add_4106_5.INIT1 = 16'h9696;
    defparam add_4106_5.INJECT1_0 = "NO";
    defparam add_4106_5.INJECT1_1 = "NO";
    CCU2C add_4106_3 (.A0(d_out_d_11__N_1888[17]), .B0(ISquare[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16756), .COUT(n16757), .S1(n90_adj_5575));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_3.INIT0 = 16'h666a;
    defparam add_4106_3.INIT1 = 16'h555f;
    defparam add_4106_3.INJECT1_0 = "NO";
    defparam add_4106_3.INJECT1_1 = "NO";
    CCU2C add_4106_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16756));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam add_4106_1.INIT0 = 16'h0000;
    defparam add_4106_1.INIT1 = 16'haaaf;
    defparam add_4106_1.INJECT1_0 = "NO";
    defparam add_4106_1.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_25 (.A0(d_tmp[58]), .B0(cout_adj_5496), .C0(n117_adj_5064), 
          .D0(n15_adj_4755), .A1(d_tmp[59]), .B1(cout_adj_5496), .C1(n114_adj_5063), 
          .D1(n14_adj_4756), .CIN(n16335), .COUT(n16336), .S0(d6_71__N_1459[58]), 
          .S1(d6_71__N_1459[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1448_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_25.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_4 (.A0(phase_inc_carrGen1[2]), .B0(phase_accum_adj_5665[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[3]), .B1(phase_accum_adj_5665[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16600), .COUT(n16601), .S0(n315), 
          .S1(n312));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_4.INIT0 = 16'h666a;
    defparam phase_accum_add_4_4.INIT1 = 16'h666a;
    defparam phase_accum_add_4_4.INJECT1_0 = "NO";
    defparam phase_accum_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_30 (.A0(d_d9_adj_5685[63]), .B0(d9_adj_5684[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[64]), .B1(d9_adj_5684[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16508), .COUT(n16509), .S0(n102_adj_4917), 
          .S1(n99_adj_4916));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_30.INJECT1_1 = "NO";
    CCU2C add_4107_65 (.A0(phase_inc_carrGen[62]), .B0(n13099), .C0(n12221), 
          .D0(n3715), .A1(phase_inc_carrGen[63]), .B1(n13099), .C1(n12223), 
          .D1(n3715), .CIN(n16750), .S0(n137), .S1(n134));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_65.INIT0 = 16'h74b8;
    defparam add_4107_65.INIT1 = 16'h74b8;
    defparam add_4107_65.INJECT1_0 = "NO";
    defparam add_4107_65.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_2 (.A0(phase_inc_carrGen1[0]), .B0(phase_accum_adj_5665[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[1]), .B1(phase_accum_adj_5665[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16600), .S1(n318));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_2.INIT0 = 16'h0008;
    defparam phase_accum_add_4_2.INIT1 = 16'h666a;
    defparam phase_accum_add_4_2.INJECT1_0 = "NO";
    defparam phase_accum_add_4_2.INJECT1_1 = "NO";
    CCU2C add_4107_63 (.A0(phase_inc_carrGen[60]), .B0(n13099), .C0(n2332), 
          .D0(n3715), .A1(phase_inc_carrGen[61]), .B1(n13099), .C1(n12219), 
          .D1(n3715), .CIN(n16749), .COUT(n16750), .S0(n143), .S1(n140));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_63.INIT0 = 16'h74b8;
    defparam add_4107_63.INIT1 = 16'h74b8;
    defparam add_4107_63.INJECT1_0 = "NO";
    defparam add_4107_63.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5663), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15392));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(62[13:22])
    defparam _add_1_1517_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1517_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1517_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_1.INJECT1_1 = "NO";
    LUT4 i5623_2_lut (.A(d2[0]), .B(d1[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5623_2_lut.init = 16'h6666;
    LUT4 i3246_2_lut_2_lut (.A(n18268), .B(n292), .Z(n2451)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i3246_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_4_lut_4_lut (.A(led_c_1), .B(led_c_0), .C(led_c_4), 
         .D(led_c_3), .Z(n17536)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_4_lut_4_lut.init = 16'h0010;
    LUT4 i5622_2_lut (.A(d3[0]), .B(d2[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5622_2_lut.init = 16'h6666;
    LUT4 mux_751_i32_3_lut (.A(led_c_2), .B(led_c_4), .C(n2845), .Z(n3716)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_751_i32_3_lut.init = 16'hc5c5;
    LUT4 i5642_2_lut (.A(d4[0]), .B(d3[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5642_2_lut.init = 16'h6666;
    LUT4 equal_300_i10_2_lut_2_lut (.A(led_c_1), .B(led_c_0), .Z(n10_adj_4574)) /* synthesis lut_function=((B)+!A) */ ;
    defparam equal_300_i10_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_326_i51_4_lut (.A(n2542), .B(n169_adj_5403), .C(n18135), 
         .D(n2593), .Z(n2342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i51_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_rep_167_3_lut_4_lut (.A(led_c_2), .B(led_c_1), .C(led_c_4), 
         .D(led_c_0), .Z(n18137)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_167_3_lut_4_lut.init = 16'h0100;
    LUT4 i3322_2_lut (.A(n163), .B(led_c_3), .Z(n2542)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3322_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_175_3_lut (.A(led_c_2), .B(led_c_1), .C(led_c_0), 
         .Z(n18145)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_175_3_lut.init = 16'h1010;
    LUT4 i5624_2_lut (.A(d1_adj_5673[0]), .B(MixerOutCos[0]), .Z(d1_71__N_418_adj_5689[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5624_2_lut.init = 16'h6666;
    LUT4 mux_751_i31_3_lut (.A(led_c_2), .B(led_c_4), .C(n2845), .Z(n3677)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_751_i31_3_lut.init = 16'h3a3a;
    LUT4 i5625_2_lut (.A(d5[0]), .B(d4[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5625_2_lut.init = 16'h6666;
    LUT4 led_c_0_bdd_3_lut (.A(led_c_1), .B(led_c_2), .C(led_c_3), .Z(n18074)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam led_c_0_bdd_3_lut.init = 16'hf6f6;
    LUT4 mux_326_i52_4_lut (.A(n12043), .B(n166_adj_5402), .C(n18135), 
         .D(n2593), .Z(n2341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i52_4_lut.init = 16'hcfca;
    VLO i1 (.Z(GND_net));
    LUT4 i2300_3_lut_4_lut (.A(n18138), .B(n18267), .C(led_c_3), .D(n211), 
         .Z(n12015)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2300_3_lut_4_lut.init = 16'hf808;
    LUT4 i6642_4_lut (.A(n17593), .B(n18142), .C(n18087), .D(n17963), 
         .Z(clk_80mhz_enable_891)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i6642_4_lut.init = 16'h3032;
    LUT4 i2292_3_lut_4_lut (.A(n18138), .B(n18267), .C(led_c_3), .D(n223), 
         .Z(n12007)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2292_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_326_i49_4_lut (.A(n10_adj_5662), .B(n175_adj_5405), .C(n18135), 
         .D(n17322), .Z(n2344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i49_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_adj_61 (.A(led_c_3), .B(n169), .Z(n10_adj_5662)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_2_lut_adj_61.init = 16'h8888;
    LUT4 i2286_3_lut_4_lut (.A(n18138), .B(led_c_2), .C(n18268), .D(n232), 
         .Z(n12001)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2286_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_326_i50_4_lut (.A(n2409), .B(n172_adj_5404), .C(n18135), 
         .D(n12136), .Z(n2343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i50_4_lut.init = 16'hcfca;
    FD1S3AX o_Rx_Byte_i3_rep_183 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(n18267));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i3_rep_183.GSR = "ENABLED";
    LUT4 i3252_2_lut (.A(n166), .B(n18268), .Z(n2409)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3252_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_179 (.A(o_Rx_DV), .B(led_c_5), .C(led_c_7), .Z(n18149)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_3_lut_rep_179.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_172_4_lut (.A(o_Rx_DV), .B(led_c_5), .C(led_c_7), 
         .D(led_c_6), .Z(n18142)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_2_lut_rep_172_4_lut.init = 16'hf7ff;
    LUT4 mux_326_i4_3_lut_4_lut (.A(led_c_3), .B(n18141), .C(n310), .D(n17322), 
         .Z(n2389)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam mux_326_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3160_rep_100_2_lut (.A(led_c_2), .B(led_c_1), .Z(n17963)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3160_rep_100_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_4_lut (.A(o_Rx_DV), .B(led_c_5), .C(led_c_7), .D(led_c_4), 
         .Z(n17319)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i1_2_lut_4_lut.init = 16'hf7ff;
    LUT4 mux_326_i2_4_lut_4_lut (.A(led_c_3), .B(n18141), .C(n18129), 
         .D(n316), .Z(n2391)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam mux_326_i2_4_lut_4_lut.init = 16'h4501;
    LUT4 mux_326_i3_4_lut_4_lut (.A(led_c_3), .B(n18141), .C(n18134), 
         .D(n313), .Z(n2390)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam mux_326_i3_4_lut_4_lut.init = 16'h4501;
    LUT4 mux_326_i47_4_lut (.A(n12035), .B(n181_adj_5407), .C(n18135), 
         .D(n2593), .Z(n2346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i47_4_lut.init = 16'hcfca;
    CCU2C add_4107_61 (.A0(phase_inc_carrGen[58]), .B0(n13099), .C0(n2334), 
          .D0(n3715), .A1(phase_inc_carrGen[59]), .B1(n13099), .C1(n2333), 
          .D1(n3715), .CIN(n16748), .COUT(n16749), .S0(n149), .S1(n146));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_61.INIT0 = 16'h74b8;
    defparam add_4107_61.INIT1 = 16'h74b8;
    defparam add_4107_61.INJECT1_0 = "NO";
    defparam add_4107_61.INJECT1_1 = "NO";
    CCU2C add_4107_59 (.A0(phase_inc_carrGen[56]), .B0(n13099), .C0(n2336), 
          .D0(n3715), .A1(phase_inc_carrGen[57]), .B1(n13099), .C1(n12217), 
          .D1(n3715), .CIN(n16747), .COUT(n16748), .S0(n155), .S1(n152));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_59.INIT0 = 16'h74b8;
    defparam add_4107_59.INIT1 = 16'h74b8;
    defparam add_4107_59.INJECT1_0 = "NO";
    defparam add_4107_59.INJECT1_1 = "NO";
    CCU2C add_4107_57 (.A0(phase_inc_carrGen[54]), .B0(n13099), .C0(n2338), 
          .D0(n3715), .A1(phase_inc_carrGen[55]), .B1(n13099), .C1(n2337), 
          .D1(n3715), .CIN(n16746), .COUT(n16747), .S0(n161), .S1(n158));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_57.INIT0 = 16'h74b8;
    defparam add_4107_57.INIT1 = 16'h74b8;
    defparam add_4107_57.INJECT1_0 = "NO";
    defparam add_4107_57.INJECT1_1 = "NO";
    CCU2C add_4107_55 (.A0(phase_inc_carrGen[52]), .B0(n13099), .C0(n12215), 
          .D0(n3715), .A1(phase_inc_carrGen[53]), .B1(n13099), .C1(n2339), 
          .D1(n3715), .CIN(n16745), .COUT(n16746), .S0(n167), .S1(n164));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_55.INIT0 = 16'h74b8;
    defparam add_4107_55.INIT1 = 16'h74b8;
    defparam add_4107_55.INJECT1_0 = "NO";
    defparam add_4107_55.INJECT1_1 = "NO";
    LUT4 i2328_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(n18268), .D(n160), 
         .Z(n12043)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2328_3_lut_4_lut.init = 16'hf404;
    \CIC(width=72,decimation_ratio=4096)  CIC1Sin (.d_tmp({d_tmp}), .clk_80mhz(clk_80mhz), 
            .d5({d5}), .d_d_tmp({d_d_tmp}), .d2({d2}), .d2_71__N_490({d2_71__N_490}), 
            .d3({d3}), .d3_71__N_562({d3_71__N_562}), .d4({d4}), .d4_71__N_634({d4_71__N_634}), 
            .d5_71__N_706({d5_71__N_706}), .d6({d6}), .d6_71__N_1459({d6_71__N_1459}), 
            .d_d6({d_d6}), .CIC1_out_clkSin(CIC1_out_clkSin), .d7({d7}), 
            .d7_71__N_1531({d7_71__N_1531}), .d_d7({d_d7}), .d8({d8}), 
            .d8_71__N_1603({d8_71__N_1603}), .d_d8({d_d8}), .d9({d9}), 
            .d9_71__N_1675({d9_71__N_1675}), .d_d9({d_d9}), .CIC1_outSin({CIC1_outSin}), 
            .d1({d1}), .d1_71__N_418({d1_71__N_418}), .count({count}), 
            .n32(n32_adj_4702), .n25(n25_adj_4709), .n24(n24_adj_4710), 
            .\CICGain[1] (CICGain[1]), .\CICGain[0] (CICGain[0]), .n9(n9_adj_4761), 
            .n8(n8_adj_4762), .n33(n33_adj_4774), .n27(n27_adj_4707), 
            .n26(n26_adj_4708), .n26_adj_115(n26_adj_4781), .n32_adj_116(n32_adj_4775), 
            .n29(n29_adj_4778), .n35(n35_adj_4810), .n35_adj_117(n35_adj_4772), 
            .\d10[69] (d10_adj_5686[69]), .\d10[68] (d10_adj_5686[68]), 
            .n34(n34_adj_4793), .\d10[65] (d10_adj_5686[65]), .\d10[66] (d10_adj_5686[66]), 
            .\d10[67] (d10_adj_5686[67]), .n11(n11_adj_4592), .n10(n10_adj_4617), 
            .n37(n37_adj_4688), .n36(n36_adj_4693), .n28(n28_adj_4779), 
            .\d10[70] (d10_adj_5686[70]), .\d10[71] (d10_adj_5686[71]), 
            .n37_adj_118(n37_adj_4812), .n34_adj_119(n34_adj_4773), .n37_adj_120(n37_adj_4770), 
            .n33_adj_121(n33_adj_4794), .n32_adj_122(n32_adj_4795), .n36_adj_123(n36_adj_4771), 
            .n31(n31_adj_4776), .n30(n30_adj_4777), .n87_adj_228({n36_adj_5090, 
            n39, n42, n45, n48, n51, n54, n57, n60, n63_adj_5091, 
            n66_adj_5092, n69, n72, n75, n78_adj_5093, n81_adj_5094}), 
            .n63_adj_125(n63), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_5711[2]), 
            .n5(n5_adj_4689), .n11_adj_126(n11_adj_4759), .n10_adj_127(n10_adj_4760), 
            .n13(n13_adj_4757), .n12(n12_adj_4758), .n15(n15_adj_4755), 
            .n4(n4_adj_4690), .n14(n14_adj_4756), .n17(n17_adj_4732), 
            .n16(n16_adj_4731), .n25_adj_128(n25_adj_4802), .n24_adj_129(n24_adj_4803), 
            .n29_adj_130(n29_adj_4705), .n28_adj_131(n28_adj_4706), .n31_adj_132(n31_adj_4703), 
            .n30_adj_133(n30_adj_4704), .n64(n64), .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_5711[3]), 
            .n36_adj_134(n36_adj_4811), .n65(n65), .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_5711[4]), 
            .n66_adj_135(n66), .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_5711[5]), 
            .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_5711[6]), .n13_adj_136(n13_adj_4576), 
            .n12_adj_137(n12_adj_4577), .\d10[64] (d10_adj_5686[64]), .n15_adj_138(n15_adj_4573), 
            .\d10[62] (d10_adj_5686[62]), .\d10[63] (d10_adj_5686[63]), 
            .n17784(n17784), .\d10[60] (d10_adj_5686[60]), .n14_adj_139(n14_adj_4575), 
            .n17_adj_140(n17_adj_4571), .\d10[61] (d10_adj_5686[61]), .n17805(n17805), 
            .\d10[59] (d10_adj_5686[59]), .n16_adj_141(n16_adj_4572), .n3(n3_adj_4767), 
            .n2(n2_adj_4768), .n19(n19_adj_4808), .n5_adj_142(n5_adj_4765), 
            .n4_adj_143(n4_adj_4766), .n7(n7_adj_4763), .n6(n6_adj_4764), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_5711[7]), .n33_adj_144(n33_adj_4701), 
            .n22(n22_adj_4836), .n6_adj_145(n6_adj_4687), .n19_adj_146(n19_adj_4569), 
            .n27_adj_147(n27), .n26_adj_148(n26), .n29_adj_149(n29), .n18(n18_adj_4570), 
            .n23(n23_adj_4804), .n22_adj_150(n22_adj_4805), .n28_adj_151(n28), 
            .n21(n21_adj_4567), .n20(n20_adj_4568), .n18_adj_152(n18_adj_4809), 
            .n31_adj_153(n31_adj_4813), .n35_adj_154(n35_adj_4699), .n34_adj_155(n34_adj_4700), 
            .n30_adj_156(n30), .n33_adj_157(n33_adj_4696), .n25_adj_158(n25), 
            .n118(n118), .n120(n120_adj_5049), .cout(cout_adj_5612), .n32_adj_159(n32_adj_4792), 
            .n24_adj_160(n24), .n115(n115), .n117(n117_adj_5048), .n35_adj_161(n35_adj_4694), 
            .n27_adj_162(n27_adj_4800), .n34_adj_163(n34_adj_4695), .n26_adj_164(n26_adj_4801), 
            .n29_adj_165(n29_adj_4798), .n112(n112), .n114(n114_adj_5047), 
            .n3_adj_166(n3_adj_4691), .n109(n109), .n111(n111_adj_5046), 
            .n106(n106), .n108(n108_adj_5045), .n103(n103), .n105(n105_adj_5044), 
            .n37_adj_167(n37_adj_4697), .n28_adj_168(n28_adj_4799), .n100(n100), 
            .n102(n102_adj_5043), .n97(n97), .n99(n99_adj_5042), .n36_adj_169(n36_adj_4698), 
            .n94(n94), .n96(n96_adj_5041), .n91(n91), .n93(n93_adj_5040), 
            .n88(n88), .n90(n90_adj_5039), .n2_adj_170(n2_adj_4692), .n85(n85), 
            .n87(n87_adj_5038), .n3_adj_171(n3_adj_4565), .n2_adj_172(n2_adj_4566), 
            .n5_adj_173(n5_adj_4729), .n4_adj_174(n4_adj_4730), .n7_adj_175(n7_adj_4727), 
            .n82(n82), .n84(n84_adj_5037), .n6_adj_176(n6_adj_4728), .n9_adj_177(n9_adj_4725), 
            .n3_adj_178(n3_adj_4834), .n8_adj_179(n8_adj_4726), .n23_adj_180(n23), 
            .n7_adj_181(n7_adj_4658), .n2_adj_182(n2_adj_4835), .n5_adj_183(n5_adj_4832), 
            .n79(n79), .n81_adj_184(n81_adj_5036), .n9_adj_185(n9_adj_4625), 
            .n76(n76), .n78_adj_186(n78_adj_5035), .n4_adj_187(n4_adj_4833), 
            .n11_adj_188(n11_adj_4723), .n10_adj_189(n10_adj_4724), .n7_adj_190(n7_adj_4830), 
            .n6_adj_191(n6_adj_4831), .n31_adj_192(n31_adj_4796), .n9_adj_193(n9_adj_4828), 
            .n21_adj_194(n21_adj_4806), .n20_adj_195(n20_adj_4807), .n8_adj_196(n8_adj_4829), 
            .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5711[10]), .n11_adj_197(n11_adj_4826), 
            .n13_adj_198(n13_adj_4721), .n12_adj_199(n12_adj_4722), .n30_adj_200(n30_adj_4797), 
            .n10_adj_201(n10_adj_4827), .n13_adj_202(n13_adj_4824), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5711[11]), 
            .n8_adj_203(n8_adj_4655), .n12_adj_204(n12_adj_4825), .n15_adj_205(n15_adj_4822), 
            .n15_adj_206(n15_adj_4719), .n14_adj_207(n14_adj_4720), .n14_adj_208(n14_adj_4823), 
            .n17_adj_209(n17_adj_4820), .n16_adj_210(n16_adj_4821), .n19_adj_211(n19_adj_4818), 
            .n17_adj_212(n17_adj_4717), .n18_adj_213(n18_adj_4819), .n16_adj_214(n16_adj_4718), 
            .n21_adj_215(n21_adj_4816), .n20_adj_216(n20_adj_4817), .n19_adj_217(n19_adj_4715), 
            .n23_adj_218(n23_adj_4814), .n22_adj_219(n22_adj_4815), .n25_adj_220(n25_adj_4782), 
            .n18_adj_221(n18_adj_4716), .n21_adj_222(n21_adj_4713), .n20_adj_223(n20_adj_4714), 
            .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_5711[8]), .n24_adj_224(n24_adj_4783), 
            .n27_adj_225(n27_adj_4780), .n23_adj_226(n23_adj_4711), .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_5711[9]), 
            .n22_adj_227(n22_adj_4712)) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(181[45] 187[2])
    LUT4 mux_326_i48_4_lut (.A(n12037), .B(n178_adj_5406), .C(n18135), 
         .D(n2593), .Z(n2345)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i48_4_lut.init = 16'hc0ca;
    LUT4 i2318_3_lut_4_lut (.A(n18267), .B(n18138), .C(n18268), .D(n178), 
         .Z(n12033)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2318_3_lut_4_lut.init = 16'hf404;
    LUT4 i5563_2_lut_rep_180 (.A(ISquare[23]), .B(ISquare[22]), .Z(n18150)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam i5563_2_lut_rep_180.init = 16'heeee;
    LUT4 mux_326_i45_4_lut (.A(n2414), .B(n187_adj_5409), .C(n18135), 
         .D(n12136), .Z(n2348)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i45_4_lut.init = 16'hc0ca;
    LUT4 i5607_1_lut_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n40)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam i5607_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i2308_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(n18268), .D(n199), 
         .Z(n12023)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2308_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_326_i46_4_lut (.A(n12033), .B(n184_adj_5408), .C(n18135), 
         .D(n2593), .Z(n2347)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i46_4_lut.init = 16'hc0ca;
    LUT4 PWMOut_I_0_1_lut (.A(PWMOutP4_c), .Z(PWMOutN4_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(139[19:26])
    defparam PWMOut_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_173_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n18143)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam i1_2_lut_rep_173_3_lut.init = 16'hfefe;
    SinCos SinCos1 (.clk_80mhz(clk_80mhz), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    LUT4 mux_326_i21_4_lut (.A(n11989), .B(n259_adj_5433), .C(n18135), 
         .D(n2593), .Z(n2372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i21_4_lut.init = 16'hcfca;
    LUT4 i2478_4_lut (.A(n262_adj_5434), .B(n256), .C(led_c_3), .D(n18141), 
         .Z(n12209)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2478_4_lut.init = 16'hcac0;
    LUT4 mux_751_i23_3_lut_rep_166 (.A(led_c_2), .B(led_c_4), .C(n2845), 
         .Z(n18136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_751_i23_3_lut_rep_166.init = 16'hcaca;
    LUT4 i2310_3_lut_4_lut (.A(n18267), .B(n18138), .C(led_c_3), .D(n196), 
         .Z(n12025)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2310_3_lut_4_lut.init = 16'hf404;
    LUT4 i2480_4_lut (.A(n256_adj_5432), .B(n250), .C(led_c_3), .D(n18141), 
         .Z(n12211)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2480_4_lut.init = 16'hcac0;
    LUT4 mux_326_i19_4_lut (.A(n11985), .B(n265_adj_5435), .C(n18135), 
         .D(n2593), .Z(n2374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i19_4_lut.init = 16'hcfca;
    PLL PLL1 (.clk_25mhz_c(clk_25mhz_c), .clk_80mhz(clk_80mhz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(145[5] 148[2])
    CCU2C _add_1_1577_add_4_12 (.A0(d4_adj_5676[45]), .B0(d3_adj_5675[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[46]), .B1(d3_adj_5675[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16272), .COUT(n16273), .S0(n156_adj_4560), 
          .S1(n153_adj_4561));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_12.INJECT1_1 = "NO";
    CCU2C add_4107_53 (.A0(phase_inc_carrGen[50]), .B0(n13099), .C0(n2342), 
          .D0(n3677), .A1(phase_inc_carrGen[51]), .B1(n13099), .C1(n2341), 
          .D1(n3715), .CIN(n16744), .COUT(n16745), .S0(n173), .S1(n170));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_53.INIT0 = 16'h74b8;
    defparam add_4107_53.INIT1 = 16'h74b8;
    defparam add_4107_53.INJECT1_0 = "NO";
    defparam add_4107_53.INJECT1_1 = "NO";
    CCU2C add_4107_51 (.A0(phase_inc_carrGen[48]), .B0(n13099), .C0(n2344), 
          .D0(n3677), .A1(phase_inc_carrGen[49]), .B1(n13099), .C1(n2343), 
          .D1(n3677), .CIN(n16743), .COUT(n16744), .S0(n179), .S1(n176));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_51.INIT0 = 16'h74b8;
    defparam add_4107_51.INIT1 = 16'h74b8;
    defparam add_4107_51.INJECT1_0 = "NO";
    defparam add_4107_51.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_17 (.A0(d4_adj_5676[50]), .B0(cout_adj_5150), 
          .C0(n141_adj_4858), .D0(d5_adj_5677[50]), .A1(d4_adj_5676[51]), 
          .B1(cout_adj_5150), .C1(n138_adj_4857), .D1(d5_adj_5677[51]), 
          .CIN(n16353), .COUT(n16354), .S0(d5_71__N_706_adj_5693[50]), 
          .S1(d5_71__N_706_adj_5693[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_17.INJECT1_1 = "NO";
    CCU2C add_4107_49 (.A0(phase_inc_carrGen[46]), .B0(n13099), .C0(n2346), 
          .D0(n11716), .A1(phase_inc_carrGen[47]), .B1(n13099), .C1(n2345), 
          .D1(n11716), .CIN(n16742), .COUT(n16743), .S0(n185), .S1(n182));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_49.INIT0 = 16'h74b8;
    defparam add_4107_49.INIT1 = 16'h74b8;
    defparam add_4107_49.INJECT1_0 = "NO";
    defparam add_4107_49.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_28 (.A0(d_d9_adj_5685[61]), .B0(d9_adj_5684[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[62]), .B1(d9_adj_5684[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16507), .COUT(n16508), .S0(n108_adj_4919), 
          .S1(n105_adj_4918));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_37 (.A0(d6[70]), .B0(cout_adj_5490), .C0(n81_adj_4961), 
          .D0(n3_adj_4565), .A1(d6[71]), .B1(cout_adj_5490), .C1(n78_adj_4960), 
          .D1(n2_adj_4566), .CIN(n16533), .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_38 (.A0(d5[71]), .B0(d4[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16598), .S0(n78_adj_5448));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1565_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_36 (.A0(d5[69]), .B0(d4[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[70]), .B1(d4[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16597), .COUT(n16598), .S0(n84_adj_5450), .S1(n81_adj_5449));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_26 (.A0(d_d9_adj_5685[59]), .B0(d9_adj_5684[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[60]), .B1(d9_adj_5684[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16506), .COUT(n16507), .S0(n114_adj_4921), 
          .S1(n111_adj_4920));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_26.INJECT1_1 = "NO";
    CCU2C add_4107_47 (.A0(phase_inc_carrGen[44]), .B0(n13099), .C0(n2348), 
          .D0(n18136), .A1(phase_inc_carrGen[45]), .B1(n13099), .C1(n2347), 
          .D1(n3715), .CIN(n16741), .COUT(n16742), .S0(n191), .S1(n188));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_47.INIT0 = 16'h74b8;
    defparam add_4107_47.INIT1 = 16'h74b8;
    defparam add_4107_47.INJECT1_0 = "NO";
    defparam add_4107_47.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_35 (.A0(d6[68]), .B0(cout_adj_5490), .C0(n87_adj_4963), 
          .D0(n5_adj_4729), .A1(d6[69]), .B1(cout_adj_5490), .C1(n84_adj_4962), 
          .D1(n4_adj_4730), .CIN(n16532), .COUT(n16533), .S0(d7_71__N_1531[68]), 
          .S1(d7_71__N_1531[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_34 (.A0(d5[67]), .B0(d4[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[68]), .B1(d4[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16596), .COUT(n16597), .S0(n90_adj_5452), .S1(n87_adj_5451));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_34.INJECT1_1 = "NO";
    LUT4 mux_326_i43_4_lut (.A(n12029), .B(n193_adj_5411), .C(n18135), 
         .D(n2593), .Z(n2350)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i43_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1565_add_4_32 (.A0(d5[65]), .B0(d4[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[66]), .B1(d4[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16595), .COUT(n16596), .S0(n96_adj_5454), .S1(n93_adj_5453));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_30 (.A0(d5[63]), .B0(d4[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[64]), .B1(d4[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16594), .COUT(n16595), .S0(n102_adj_5456), .S1(n99_adj_5455));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_28 (.A0(d5[61]), .B0(d4[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[62]), .B1(d4[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16593), .COUT(n16594), .S0(n108_adj_5458), .S1(n105_adj_5457));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_26 (.A0(d5[59]), .B0(d4[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[60]), .B1(d4[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16592), .COUT(n16593), .S0(n114_adj_5460), .S1(n111_adj_5459));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_24 (.A0(d5[57]), .B0(d4[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[58]), .B1(d4[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16591), .COUT(n16592), .S0(n120_adj_5462), .S1(n117_adj_5461));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_24.INJECT1_1 = "NO";
    LUT4 i2006_1_lut_3_lut (.A(led_c_2), .B(led_c_4), .C(n2845), .Z(n11716)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2006_1_lut_3_lut.init = 16'h3535;
    CCU2C _add_1_1565_add_4_22 (.A0(d5[55]), .B0(d4[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[56]), .B1(d4[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16590), .COUT(n16591), .S0(n126_adj_5464), .S1(n123_adj_5463));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_35 (.A0(d4_adj_5676[68]), .B0(cout_adj_5150), 
          .C0(n87_adj_4840), .D0(d5_adj_5677[68]), .A1(d4_adj_5676[69]), 
          .B1(cout_adj_5150), .C1(n84_adj_4839), .D1(d5_adj_5677[69]), 
          .CIN(n16362), .COUT(n16363), .S0(d5_71__N_706_adj_5693[68]), 
          .S1(d5_71__N_706_adj_5693[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_20 (.A0(d5[53]), .B0(d4[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[54]), .B1(d4[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16589), .COUT(n16590), .S0(n132_adj_5466), .S1(n129_adj_5465));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_18 (.A0(d5[51]), .B0(d4[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[52]), .B1(d4[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16588), .COUT(n16589), .S0(n138_adj_5468), .S1(n135_adj_5467));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_18.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i1 (.D(o_Rx_Byte1[0]), .CK(clk_80mhz), .Q(led_c_0));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    CCU2C _add_1_1637_add_4_24 (.A0(d_d9_adj_5685[57]), .B0(d9_adj_5684[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[58]), .B1(d9_adj_5684[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16505), .COUT(n16506), .S0(n120_adj_4923), 
          .S1(n117_adj_4922));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_33 (.A0(d6[66]), .B0(cout_adj_5490), .C0(n93_adj_4965), 
          .D0(n7_adj_4727), .A1(d6[67]), .B1(cout_adj_5490), .C1(n90_adj_4964), 
          .D1(n6_adj_4728), .CIN(n16531), .COUT(n16532), .S0(d7_71__N_1531[66]), 
          .S1(d7_71__N_1531[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_16 (.A0(d5[49]), .B0(d4[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[50]), .B1(d4[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16587), .COUT(n16588), .S0(n144_adj_5470), .S1(n141_adj_5469));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_16.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i4_rep_184 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(n18268));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam o_Rx_Byte_i4_rep_184.GSR = "ENABLED";
    CCU2C _add_1_1565_add_4_14 (.A0(d5[47]), .B0(d4[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[48]), .B1(d4[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16586), .COUT(n16587), .S0(n150_adj_5472), .S1(n147_adj_5471));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_12 (.A0(d5[45]), .B0(d4[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[46]), .B1(d4[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16585), .COUT(n16586), .S0(n156_adj_5474), .S1(n153_adj_5473));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_31 (.A0(d6[64]), .B0(cout_adj_5490), .C0(n99_adj_4967), 
          .D0(n9_adj_4725), .A1(d6[65]), .B1(cout_adj_5490), .C1(n96_adj_4966), 
          .D1(n8_adj_4726), .CIN(n16530), .COUT(n16531), .S0(d7_71__N_1531[64]), 
          .S1(d7_71__N_1531[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_10 (.A0(d5[43]), .B0(d4[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[44]), .B1(d4[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16584), .COUT(n16585), .S0(n162_adj_5476), .S1(n159_adj_5475));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_10.INJECT1_1 = "NO";
    CCU2C add_4107_45 (.A0(phase_inc_carrGen[42]), .B0(n13099), .C0(n2350), 
          .D0(n18131), .A1(phase_inc_carrGen[43]), .B1(n13099), .C1(n2349), 
          .D1(n3685), .CIN(n16740), .COUT(n16741), .S0(n197), .S1(n194));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_45.INIT0 = 16'h74b8;
    defparam add_4107_45.INIT1 = 16'h74b8;
    defparam add_4107_45.INJECT1_0 = "NO";
    defparam add_4107_45.INJECT1_1 = "NO";
    LUT4 i2304_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(led_c_3), .D(n205), 
         .Z(n12019)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2304_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_326_i44_4_lut (.A(n12031), .B(n190_adj_5410), .C(n18135), 
         .D(n2593), .Z(n2349)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i44_4_lut.init = 16'hc0ca;
    PFUMX i6720 (.BLUT(n18189), .ALUT(n18190), .C0(led_c_2), .Z(n18191));
    CCU2C _add_1_1577_add_4_34 (.A0(d4_adj_5676[67]), .B0(d3_adj_5675[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[68]), .B1(d3_adj_5675[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16283), .COUT(n16284), .S0(n90), 
          .S1(n87));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_30 (.A0(d4_adj_5676[63]), .B0(d3_adj_5675[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[64]), .B1(d3_adj_5675[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16281), .COUT(n16282), .S0(n102), 
          .S1(n99));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_32 (.A0(d4_adj_5676[65]), .B0(d3_adj_5675[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5676[66]), .B1(d3_adj_5675[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16282), .COUT(n16283), .S0(n96), 
          .S1(n93));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1577_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_32.INJECT1_1 = "NO";
    LUT4 i2274_3_lut_4_lut (.A(n18138), .B(n18267), .C(led_c_3), .D(n253), 
         .Z(n11989)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2274_3_lut_4_lut.init = 16'hf707;
    LUT4 i26_4_lut_adj_62 (.A(n2593), .B(n199_adj_5413), .C(n18135), .D(n13_adj_5488), 
         .Z(n11_adj_5487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i26_4_lut_adj_62.init = 16'hcacf;
    LUT4 mux_326_i17_4_lut (.A(n11981), .B(n271_adj_5437), .C(n18135), 
         .D(n2593), .Z(n2376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i17_4_lut.init = 16'hcfca;
    CCU2C _add_1_1463_add_4_29 (.A0(d6[62]), .B0(cout_adj_5490), .C0(n105_adj_4969), 
          .D0(n11_adj_4723), .A1(d6[63]), .B1(cout_adj_5490), .C1(n102_adj_4968), 
          .D1(n10_adj_4724), .CIN(n16529), .COUT(n16530), .S0(d7_71__N_1531[62]), 
          .S1(d7_71__N_1531[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_29.INJECT1_1 = "NO";
    CCU2C add_4107_43 (.A0(phase_inc_carrGen[40]), .B0(n13099), .C0(n11_adj_5487), 
          .D0(n3677), .A1(phase_inc_carrGen[41]), .B1(n13099), .C1(n12213), 
          .D1(n3685), .CIN(n16739), .COUT(n16740), .S0(n203), .S1(n200));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_43.INIT0 = 16'h74b8;
    defparam add_4107_43.INIT1 = 16'h74b8;
    defparam add_4107_43.INJECT1_0 = "NO";
    defparam add_4107_43.INJECT1_1 = "NO";
    LUT4 i2482_4_lut (.A(n196_adj_5412), .B(n190), .C(led_c_3), .D(n18141), 
         .Z(n12213)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2482_4_lut.init = 16'hcac0;
    CCU2C _add_1_1463_add_4_27 (.A0(d6[60]), .B0(cout_adj_5490), .C0(n111_adj_4971), 
          .D0(n13_adj_4721), .A1(d6[61]), .B1(cout_adj_5490), .C1(n108_adj_4970), 
          .D1(n12_adj_4722), .CIN(n16528), .COUT(n16529), .S0(d7_71__N_1531[60]), 
          .S1(d7_71__N_1531[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_27.INJECT1_1 = "NO";
    CCU2C add_4107_41 (.A0(phase_inc_carrGen[38]), .B0(n13099), .C0(n2354), 
          .D0(n3715), .A1(phase_inc_carrGen[39]), .B1(n13099), .C1(n2353), 
          .D1(n3715), .CIN(n16738), .COUT(n16739), .S0(n209_adj_4996), 
          .S1(n206));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_41.INIT0 = 16'h74b8;
    defparam add_4107_41.INIT1 = 16'h74b8;
    defparam add_4107_41.INJECT1_0 = "NO";
    defparam add_4107_41.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_25 (.A0(d6[58]), .B0(cout_adj_5490), .C0(n117_adj_4973), 
          .D0(n15_adj_4719), .A1(d6[59]), .B1(cout_adj_5490), .C1(n114_adj_4972), 
          .D1(n14_adj_4720), .CIN(n16527), .COUT(n16528), .S0(d7_71__N_1531[58]), 
          .S1(d7_71__N_1531[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_25.INJECT1_1 = "NO";
    CCU2C add_4107_39 (.A0(phase_inc_carrGen[36]), .B0(n13099), .C0(n2356), 
          .D0(n18136), .A1(phase_inc_carrGen[37]), .B1(n13099), .C1(n2355), 
          .D1(n3720), .CIN(n16737), .COUT(n16738), .S0(n215), .S1(n212));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_39.INIT0 = 16'h74b8;
    defparam add_4107_39.INIT1 = 16'h74b8;
    defparam add_4107_39.INJECT1_0 = "NO";
    defparam add_4107_39.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_23 (.A0(d6[56]), .B0(cout_adj_5490), .C0(n123_adj_4975), 
          .D0(n17_adj_4717), .A1(d6[57]), .B1(cout_adj_5490), .C1(n120_adj_4974), 
          .D1(n16_adj_4718), .CIN(n16526), .COUT(n16527), .S0(d7_71__N_1531[56]), 
          .S1(d7_71__N_1531[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_23.INJECT1_1 = "NO";
    CCU2C add_4107_37 (.A0(phase_inc_carrGen[34]), .B0(n13099), .C0(n2358), 
          .D0(n18136), .A1(phase_inc_carrGen[35]), .B1(n13099), .C1(n2357), 
          .D1(n3715), .CIN(n16736), .COUT(n16737), .S0(n221), .S1(n218));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_37.INIT0 = 16'h74b8;
    defparam add_4107_37.INIT1 = 16'h74b8;
    defparam add_4107_37.INJECT1_0 = "NO";
    defparam add_4107_37.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_21 (.A0(d6[54]), .B0(cout_adj_5490), .C0(n129_adj_4977), 
          .D0(n19_adj_4715), .A1(d6[55]), .B1(cout_adj_5490), .C1(n126_adj_4976), 
          .D1(n18_adj_4716), .CIN(n16525), .COUT(n16526), .S0(d7_71__N_1531[54]), 
          .S1(d7_71__N_1531[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_21.INJECT1_1 = "NO";
    CCU2C add_4107_35 (.A0(phase_inc_carrGen[32]), .B0(n13099), .C0(n2360), 
          .D0(n3677), .A1(phase_inc_carrGen[33]), .B1(n13099), .C1(n2359), 
          .D1(n3720), .CIN(n16735), .COUT(n16736), .S0(n227), .S1(n224));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_35.INIT0 = 16'h74b8;
    defparam add_4107_35.INIT1 = 16'h74b8;
    defparam add_4107_35.INJECT1_0 = "NO";
    defparam add_4107_35.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_19 (.A0(d6[52]), .B0(cout_adj_5490), .C0(n135_adj_4979), 
          .D0(n21_adj_4713), .A1(d6[53]), .B1(cout_adj_5490), .C1(n132_adj_4978), 
          .D1(n20_adj_4714), .CIN(n16524), .COUT(n16525), .S0(d7_71__N_1531[52]), 
          .S1(d7_71__N_1531[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_19.INJECT1_1 = "NO";
    CCU2C add_4107_33 (.A0(phase_inc_carrGen[30]), .B0(n13099), .C0(n2362), 
          .D0(n3677), .A1(phase_inc_carrGen[31]), .B1(n13099), .C1(n2361), 
          .D1(n3716), .CIN(n16734), .COUT(n16735), .S0(n233), .S1(n230));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_33.INIT0 = 16'h74b8;
    defparam add_4107_33.INIT1 = 16'h74b8;
    defparam add_4107_33.INJECT1_0 = "NO";
    defparam add_4107_33.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_17 (.A0(d6[50]), .B0(cout_adj_5490), .C0(n141_adj_4981), 
          .D0(n23_adj_4711), .A1(d6[51]), .B1(cout_adj_5490), .C1(n138_adj_4980), 
          .D1(n22_adj_4712), .CIN(n16523), .COUT(n16524), .S0(d7_71__N_1531[50]), 
          .S1(d7_71__N_1531[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_17.INJECT1_1 = "NO";
    CCU2C add_4107_31 (.A0(phase_inc_carrGen[28]), .B0(n13099), .C0(n2364), 
          .D0(n3685), .A1(phase_inc_carrGen[29]), .B1(n13099), .C1(n2363), 
          .D1(n18131), .CIN(n16733), .COUT(n16734), .S0(n239), .S1(n236));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_31.INIT0 = 16'h74b8;
    defparam add_4107_31.INIT1 = 16'h74b8;
    defparam add_4107_31.INJECT1_0 = "NO";
    defparam add_4107_31.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_15 (.A0(d6[48]), .B0(cout_adj_5490), .C0(n147_adj_4983), 
          .D0(n25_adj_4709), .A1(d6[49]), .B1(cout_adj_5490), .C1(n144_adj_4982), 
          .D1(n24_adj_4710), .CIN(n16522), .COUT(n16523), .S0(d7_71__N_1531[48]), 
          .S1(d7_71__N_1531[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_15.INJECT1_1 = "NO";
    CCU2C add_4107_29 (.A0(phase_inc_carrGen[26]), .B0(n13099), .C0(n2366), 
          .D0(n3715), .A1(phase_inc_carrGen[27]), .B1(n13099), .C1(n2365), 
          .D1(n3720), .CIN(n16732), .COUT(n16733), .S0(n245), .S1(n242));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_29.INIT0 = 16'h74b8;
    defparam add_4107_29.INIT1 = 16'h74b8;
    defparam add_4107_29.INJECT1_0 = "NO";
    defparam add_4107_29.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_13 (.A0(d6[46]), .B0(cout_adj_5490), .C0(n153_adj_4985), 
          .D0(n27_adj_4707), .A1(d6[47]), .B1(cout_adj_5490), .C1(n150_adj_4984), 
          .D1(n26_adj_4708), .CIN(n16521), .COUT(n16522), .S0(d7_71__N_1531[46]), 
          .S1(d7_71__N_1531[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_13.INJECT1_1 = "NO";
    CCU2C add_4107_27 (.A0(phase_inc_carrGen[24]), .B0(n13099), .C0(n2368), 
          .D0(n3715), .A1(phase_inc_carrGen[25]), .B1(n13099), .C1(n2367), 
          .D1(n3715), .CIN(n16731), .COUT(n16732), .S0(n251), .S1(n248));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_27.INIT0 = 16'h74b8;
    defparam add_4107_27.INIT1 = 16'h74b8;
    defparam add_4107_27.INJECT1_0 = "NO";
    defparam add_4107_27.INJECT1_1 = "NO";
    CCU2C add_4107_25 (.A0(phase_inc_carrGen[22]), .B0(n13099), .C0(n11_adj_5484), 
          .D0(n18136), .A1(phase_inc_carrGen[23]), .B1(n13099), .C1(n2369), 
          .D1(n18131), .CIN(n16730), .COUT(n16731), .S0(n257), .S1(n254));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_25.INIT0 = 16'h74b8;
    defparam add_4107_25.INIT1 = 16'h74b8;
    defparam add_4107_25.INJECT1_0 = "NO";
    defparam add_4107_25.INJECT1_1 = "NO";
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 i2302_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(n18268), .D(n208), 
         .Z(n12017)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2302_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1565_add_4_8 (.A0(d5[41]), .B0(d4[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[42]), .B1(d4[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16583), .COUT(n16584), .S0(n168_adj_5478), .S1(n165_adj_5477));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_8.INJECT1_1 = "NO";
    LUT4 mux_326_i39_4_lut (.A(n12023), .B(n205_adj_5415), .C(n18135), 
         .D(n2593), .Z(n2354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i39_4_lut.init = 16'hcfca;
    LUT4 mux_326_i40_4_lut (.A(n12025), .B(n202_adj_5414), .C(n18135), 
         .D(n2593), .Z(n2353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i40_4_lut.init = 16'hcfca;
    CCU2C _add_1_1565_add_4_6 (.A0(d5[39]), .B0(d4[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[40]), .B1(d4[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16582), .COUT(n16583), .S0(n174_adj_5480), .S1(n171_adj_5479));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_4 (.A0(d5[37]), .B0(d4[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[38]), .B1(d4[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16581), .COUT(n16582), .S0(n180_adj_5482), .S1(n177_adj_5481));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_4.INJECT1_1 = "NO";
    LUT4 mux_326_i37_4_lut (.A(n12019), .B(n211_adj_5417), .C(n18135), 
         .D(n2593), .Z(n2356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i37_4_lut.init = 16'hcfca;
    LUT4 i5591_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n15364)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam i5591_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i2254_3_lut_4_lut (.A(n18138), .B(led_c_2), .C(led_c_3), .D(n289), 
         .Z(n11969)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2254_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_326_i38_4_lut (.A(n12021), .B(n208_adj_5416), .C(n18135), 
         .D(n2593), .Z(n2355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i38_4_lut.init = 16'hcfca;
    LUT4 i3171_2_lut (.A(led_c_4), .B(n2845), .Z(n3720)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i3171_2_lut.init = 16'hbbbb;
    FD1P3AX phase_inc_carrGen_i0_i0 (.D(n323), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    LUT4 i5581_1_lut_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n49)) /* synthesis lut_function=(!(A+(B))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam i5581_1_lut_2_lut.init = 16'h1111;
    LUT4 i2294_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(n18268), .D(n220), 
         .Z(n12009)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2294_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1565_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[36]), .B1(d4[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16581), .S1(n183_adj_5483));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(70[13:20])
    defparam _add_1_1565_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1565_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_2.INJECT1_1 = "NO";
    LUT4 mux_326_i35_4_lut (.A(n12015), .B(n217_adj_5419), .C(n18135), 
         .D(n2593), .Z(n2358)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i35_4_lut.init = 16'hc0ca;
    LUT4 i3176_4_lut (.A(n10_adj_4574), .B(n17595), .C(n17310), .D(n17319), 
         .Z(n12912)) /* synthesis lut_function=(A (B+(D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i3176_4_lut.init = 16'hfac8;
    LUT4 i2288_3_lut_4_lut (.A(n18267), .B(n18138), .C(led_c_3), .D(n229), 
         .Z(n12003)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2288_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_326_i36_4_lut (.A(n12017), .B(n214_adj_5418), .C(n18135), 
         .D(n2593), .Z(n2357)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i36_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1460_add_4_13 (.A0(LOCosine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16580), .S0(MixerOutCos_11__N_250[11]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1460_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1460_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_13.INJECT1_1 = "NO";
    LUT4 i2278_3_lut_4_lut (.A(n18267), .B(n18138), .C(n18268), .D(n244), 
         .Z(n11993)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2278_3_lut_4_lut.init = 16'hf404;
    LUT4 i2256_3_lut_4_lut (.A(n18138), .B(n18267), .C(n18268), .D(n286), 
         .Z(n11971)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(248[8] 284[4])
    defparam i2256_3_lut_4_lut.init = 16'hf707;
    CCU2C _add_1_1460_add_4_11 (.A0(LOCosine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16579), .COUT(n16580), .S0(MixerOutCos_11__N_250[9]), 
          .S1(MixerOutCos_11__N_250[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1460_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1460_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_11.INJECT1_1 = "NO";
    LUT4 mux_326_i33_4_lut (.A(n12011), .B(n223_adj_5421), .C(n18135), 
         .D(n2593), .Z(n2360)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i33_4_lut.init = 16'hc0ca;
    LUT4 mux_326_i34_4_lut (.A(n12013), .B(n220_adj_5420), .C(n18135), 
         .D(n2593), .Z(n2359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i34_4_lut.init = 16'hcfca;
    CCU2C _add_1_1460_add_4_9 (.A0(LOCosine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16578), .COUT(n16579), .S0(MixerOutCos_11__N_250[7]), 
          .S1(MixerOutCos_11__N_250[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1460_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1460_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_7 (.A0(LOCosine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16577), .COUT(n16578), .S0(MixerOutCos_11__N_250[5]), 
          .S1(MixerOutCos_11__N_250[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1460_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1460_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_11 (.A0(d6[44]), .B0(cout_adj_5490), .C0(n159_adj_4987), 
          .D0(n29_adj_4705), .A1(d6[45]), .B1(cout_adj_5490), .C1(n156_adj_4986), 
          .D1(n28_adj_4706), .CIN(n16520), .COUT(n16521), .S0(d7_71__N_1531[44]), 
          .S1(d7_71__N_1531[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_5 (.A0(LOCosine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16576), .COUT(n16577), .S0(MixerOutCos_11__N_250[3]), 
          .S1(MixerOutCos_11__N_250[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1460_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1460_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_3 (.A0(LOCosine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16575), .COUT(n16576), .S0(MixerOutCos_11__N_250[1]), 
          .S1(MixerOutCos_11__N_250[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1460_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1460_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16575), .S1(MixerOutCos_11__N_250[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(42[26:33])
    defparam _add_1_1460_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1460_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1460_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_1.INJECT1_1 = "NO";
    LUT4 equal_299_i11_2_lut (.A(led_c_2), .B(n18268), .Z(n11_adj_4564)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_299_i11_2_lut.init = 16'heeee;
    CCU2C _add_1_1637_add_4_22 (.A0(d_d9_adj_5685[55]), .B0(d9_adj_5684[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[56]), .B1(d9_adj_5684[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16504), .COUT(n16505));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_9 (.A0(d6[42]), .B0(cout_adj_5490), .C0(n165_adj_4989), 
          .D0(n31_adj_4703), .A1(d6[43]), .B1(cout_adj_5490), .C1(n162_adj_4988), 
          .D1(n30_adj_4704), .CIN(n16519), .COUT(n16520), .S0(d7_71__N_1531[42]), 
          .S1(d7_71__N_1531[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_37 (.A0(d6_adj_5678[70]), .B0(cout_adj_5192), 
          .C0(n81_adj_5355), .D0(n3), .A1(d6_adj_5678[71]), .B1(cout_adj_5192), 
          .C1(n78_adj_5354), .D1(n2), .CIN(n16573), .S0(d7_71__N_1531_adj_5706[70]), 
          .S1(d7_71__N_1531_adj_5706[71]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_35 (.A0(d6_adj_5678[68]), .B0(cout_adj_5192), 
          .C0(n87_adj_5357), .D0(n5), .A1(d6_adj_5678[69]), .B1(cout_adj_5192), 
          .C1(n84_adj_5356), .D1(n4), .CIN(n16572), .COUT(n16573), .S0(d7_71__N_1531_adj_5706[68]), 
          .S1(d7_71__N_1531_adj_5706[69]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_33 (.A0(d6_adj_5678[66]), .B0(cout_adj_5192), 
          .C0(n93_adj_5359), .D0(n7), .A1(d6_adj_5678[67]), .B1(cout_adj_5192), 
          .C1(n90_adj_5358), .D1(n6), .CIN(n16571), .COUT(n16572), .S0(d7_71__N_1531_adj_5706[66]), 
          .S1(d7_71__N_1531_adj_5706[67]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_31 (.A0(d6_adj_5678[64]), .B0(cout_adj_5192), 
          .C0(n99_adj_5361), .D0(n9_adj_4682), .A1(d6_adj_5678[65]), .B1(cout_adj_5192), 
          .C1(n96_adj_5360), .D1(n8_adj_4686), .CIN(n16570), .COUT(n16571), 
          .S0(d7_71__N_1531_adj_5706[64]), .S1(d7_71__N_1531_adj_5706[65]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_31.INJECT1_1 = "NO";
    LUT4 i2266_3_lut_4_lut (.A(led_c_2), .B(n18138), .C(led_c_3), .D(n265), 
         .Z(n11981)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2266_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_326_i31_4_lut (.A(n12007), .B(n229_adj_5423), .C(n18135), 
         .D(n2593), .Z(n2362)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i31_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_174_3_lut (.A(led_c_1), .B(led_c_4), .C(led_c_0), 
         .Z(n18144)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_rep_174_3_lut.init = 16'h0202;
    nco_sig ncoGen (.\phase_accum[63] (phase_accum[63]), .sinGen_c(sinGen_c)) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(161[10] 167[2])
    CCU2C _add_1_1478_add_4_29 (.A0(d6_adj_5678[62]), .B0(cout_adj_5192), 
          .C0(n105_adj_5363), .D0(n11_adj_4684), .A1(d6_adj_5678[63]), 
          .B1(cout_adj_5192), .C1(n102_adj_5362), .D1(n10_adj_4683), .CIN(n16569), 
          .COUT(n16570), .S0(d7_71__N_1531_adj_5706[62]), .S1(d7_71__N_1531_adj_5706[63]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_27 (.A0(d6_adj_5678[60]), .B0(cout_adj_5192), 
          .C0(n111_adj_5365), .D0(n13_adj_4681), .A1(d6_adj_5678[61]), 
          .B1(cout_adj_5192), .C1(n108_adj_5364), .D1(n12_adj_4685), .CIN(n16568), 
          .COUT(n16569), .S0(d7_71__N_1531_adj_5706[60]), .S1(d7_71__N_1531_adj_5706[61]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_20 (.A0(d_d9_adj_5685[53]), .B0(d9_adj_5684[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[54]), .B1(d9_adj_5684[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16503), .COUT(n16504));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_7 (.A0(d6[40]), .B0(cout_adj_5490), .C0(n171_adj_4991), 
          .D0(n33_adj_4701), .A1(d6[41]), .B1(cout_adj_5490), .C1(n168_adj_4990), 
          .D1(n32_adj_4702), .CIN(n16518), .COUT(n16519), .S0(d7_71__N_1531[40]), 
          .S1(d7_71__N_1531[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_25 (.A0(d6_adj_5678[58]), .B0(cout_adj_5192), 
          .C0(n117_adj_5367), .D0(n15_adj_4679), .A1(d6_adj_5678[59]), 
          .B1(cout_adj_5192), .C1(n114_adj_5366), .D1(n14_adj_4680), .CIN(n16567), 
          .COUT(n16568), .S0(d7_71__N_1531_adj_5706[58]), .S1(d7_71__N_1531_adj_5706[59]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_23 (.A0(d6_adj_5678[56]), .B0(cout_adj_5192), 
          .C0(n123_adj_5369), .D0(n17_adj_4677), .A1(d6_adj_5678[57]), 
          .B1(cout_adj_5192), .C1(n120_adj_5368), .D1(n16_adj_4678), .CIN(n16566), 
          .COUT(n16567), .S0(d7_71__N_1531_adj_5706[56]), .S1(d7_71__N_1531_adj_5706[57]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_21 (.A0(d6_adj_5678[54]), .B0(cout_adj_5192), 
          .C0(n129_adj_5371), .D0(n19_adj_4675), .A1(d6_adj_5678[55]), 
          .B1(cout_adj_5192), .C1(n126_adj_5370), .D1(n18_adj_4676), .CIN(n16565), 
          .COUT(n16566), .S0(d7_71__N_1531_adj_5706[54]), .S1(d7_71__N_1531_adj_5706[55]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_19 (.A0(d6_adj_5678[52]), .B0(cout_adj_5192), 
          .C0(n135_adj_5373), .D0(n21_adj_4673), .A1(d6_adj_5678[53]), 
          .B1(cout_adj_5192), .C1(n132_adj_5372), .D1(n20_adj_4674), .CIN(n16564), 
          .COUT(n16565), .S0(d7_71__N_1531_adj_5706[52]), .S1(d7_71__N_1531_adj_5706[53]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_17 (.A0(d6_adj_5678[50]), .B0(cout_adj_5192), 
          .C0(n141_adj_5375), .D0(n23_adj_4671), .A1(d6_adj_5678[51]), 
          .B1(cout_adj_5192), .C1(n138_adj_5374), .D1(n22_adj_4672), .CIN(n16563), 
          .COUT(n16564), .S0(d7_71__N_1531_adj_5706[50]), .S1(d7_71__N_1531_adj_5706[51]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_15 (.A0(d6_adj_5678[48]), .B0(cout_adj_5192), 
          .C0(n147_adj_5377), .D0(n25_adj_4669), .A1(d6_adj_5678[49]), 
          .B1(cout_adj_5192), .C1(n144_adj_5376), .D1(n24_adj_4670), .CIN(n16562), 
          .COUT(n16563), .S0(d7_71__N_1531_adj_5706[48]), .S1(d7_71__N_1531_adj_5706[49]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_13 (.A0(d6_adj_5678[46]), .B0(cout_adj_5192), 
          .C0(n153_adj_5379), .D0(n27_adj_4667), .A1(d6_adj_5678[47]), 
          .B1(cout_adj_5192), .C1(n150_adj_5378), .D1(n26_adj_4668), .CIN(n16561), 
          .COUT(n16562), .S0(d7_71__N_1531_adj_5706[46]), .S1(d7_71__N_1531_adj_5706[47]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_11 (.A0(d6_adj_5678[44]), .B0(cout_adj_5192), 
          .C0(n159_adj_5381), .D0(n29_adj_4665), .A1(d6_adj_5678[45]), 
          .B1(cout_adj_5192), .C1(n156_adj_5380), .D1(n28_adj_4666), .CIN(n16560), 
          .COUT(n16561), .S0(d7_71__N_1531_adj_5706[44]), .S1(d7_71__N_1531_adj_5706[45]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_9 (.A0(d6_adj_5678[42]), .B0(cout_adj_5192), 
          .C0(n165_adj_5383), .D0(n31_adj_4663), .A1(d6_adj_5678[43]), 
          .B1(cout_adj_5192), .C1(n162_adj_5382), .D1(n30_adj_4664), .CIN(n16559), 
          .COUT(n16560), .S0(d7_71__N_1531_adj_5706[42]), .S1(d7_71__N_1531_adj_5706[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_5 (.A0(d6[38]), .B0(cout_adj_5490), .C0(n177_adj_4993), 
          .D0(n35_adj_4699), .A1(d6[39]), .B1(cout_adj_5490), .C1(n174_adj_4992), 
          .D1(n34_adj_4700), .CIN(n16517), .COUT(n16518), .S0(d7_71__N_1531[38]), 
          .S1(d7_71__N_1531[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_7 (.A0(d6_adj_5678[40]), .B0(cout_adj_5192), 
          .C0(n171_adj_5385), .D0(n33_adj_4661), .A1(d6_adj_5678[41]), 
          .B1(cout_adj_5192), .C1(n168_adj_5384), .D1(n32_adj_4662), .CIN(n16558), 
          .COUT(n16559), .S0(d7_71__N_1531_adj_5706[40]), .S1(d7_71__N_1531_adj_5706[41]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_7.INJECT1_1 = "NO";
    LUT4 i2258_3_lut_4_lut (.A(n18267), .B(n18138), .C(led_c_3), .D(n283), 
         .Z(n11973)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam i2258_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1637_add_4_18 (.A0(d_d9_adj_5685[51]), .B0(d9_adj_5684[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[52]), .B1(d9_adj_5684[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16502), .COUT(n16503));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_3 (.A0(d6[36]), .B0(cout_adj_5490), .C0(n183_adj_4995), 
          .D0(n37_adj_4697), .A1(d6[37]), .B1(cout_adj_5490), .C1(n180_adj_4994), 
          .D1(n36_adj_4698), .CIN(n16516), .COUT(n16517), .S0(d7_71__N_1531[36]), 
          .S1(d7_71__N_1531[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_5 (.A0(d6_adj_5678[38]), .B0(cout_adj_5192), 
          .C0(n177_adj_5387), .D0(n35_adj_4659), .A1(d6_adj_5678[39]), 
          .B1(cout_adj_5192), .C1(n174_adj_5386), .D1(n34_adj_4660), .CIN(n16557), 
          .COUT(n16558), .S0(d7_71__N_1531_adj_5706[38]), .S1(d7_71__N_1531_adj_5706[39]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_9 (.A0(d_tmp_adj_5671[42]), .B0(cout_adj_5489), 
          .C0(n165_adj_5347), .D0(n31), .A1(d_tmp_adj_5671[43]), .B1(cout_adj_5489), 
          .C1(n162_adj_5346), .D1(n30_adj_2748), .CIN(n16460), .COUT(n16461), 
          .S0(d6_71__N_1459_adj_5705[42]), .S1(d6_71__N_1459_adj_5705[43]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5490), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16516));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1463_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1463_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_3 (.A0(d6_adj_5678[36]), .B0(cout_adj_5192), 
          .C0(n183_adj_5389), .D0(n37_adj_4656), .A1(d6_adj_5678[37]), 
          .B1(cout_adj_5192), .C1(n180_adj_5388), .D1(n36_adj_4657), .CIN(n16556), 
          .COUT(n16557), .S0(d7_71__N_1531_adj_5706[36]), .S1(d7_71__N_1531_adj_5706[37]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5192), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16556));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1478_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1478_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_1.INJECT1_1 = "NO";
    CCU2C add_4107_23 (.A0(phase_inc_carrGen[20]), .B0(n13099), .C0(n2372), 
          .D0(n3715), .A1(phase_inc_carrGen[21]), .B1(n13099), .C1(n12211), 
          .D1(n3677), .CIN(n16729), .COUT(n16730), .S0(n263), .S1(n260));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_23.INIT0 = 16'h74b8;
    defparam add_4107_23.INIT1 = 16'h74b8;
    defparam add_4107_23.INJECT1_0 = "NO";
    defparam add_4107_23.INJECT1_1 = "NO";
    LUT4 mux_326_i32_4_lut (.A(n12009), .B(n226_adj_5422), .C(n18135), 
         .D(n2593), .Z(n2361)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam mux_326_i32_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1562_add_4_38 (.A0(d4[71]), .B0(d3[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16552), .S0(n78_adj_5267));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1562_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_38.INJECT1_1 = "NO";
    CCU2C add_4107_21 (.A0(phase_inc_carrGen[18]), .B0(n13099), .C0(n2374), 
          .D0(n18131), .A1(phase_inc_carrGen[19]), .B1(n13099), .C1(n12209), 
          .D1(n3720), .CIN(n16728), .COUT(n16729), .S0(n269), .S1(n266));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_21.INIT0 = 16'h74b8;
    defparam add_4107_21.INIT1 = 16'h74b8;
    defparam add_4107_21.INJECT1_0 = "NO";
    defparam add_4107_21.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_36 (.A0(d4[69]), .B0(d3[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[70]), .B1(d3[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16551), .COUT(n16552), .S0(n84_adj_5269), .S1(n81_adj_5268));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_34 (.A0(d4[67]), .B0(d3[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[68]), .B1(d3[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16550), .COUT(n16551), .S0(n90_adj_5271), .S1(n87_adj_5270));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_32 (.A0(d4[65]), .B0(d3[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[66]), .B1(d3[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16549), .COUT(n16550), .S0(n96_adj_5273), .S1(n93_adj_5272));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_32.INJECT1_1 = "NO";
    CCU2C add_4107_19 (.A0(phase_inc_carrGen[16]), .B0(n13099), .C0(n2376), 
          .D0(n3716), .A1(phase_inc_carrGen[17]), .B1(n13099), .C1(n2375), 
          .D1(n11716), .CIN(n16727), .COUT(n16728), .S0(n275), .S1(n272));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_19.INIT0 = 16'h74b8;
    defparam add_4107_19.INIT1 = 16'h74b8;
    defparam add_4107_19.INJECT1_0 = "NO";
    defparam add_4107_19.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_38 (.A0(d_d9_adj_5685[71]), .B0(d9_adj_5684[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16512), .S0(n78_adj_4909));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1637_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_30 (.A0(d4[63]), .B0(d3[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[64]), .B1(d3[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16548), .COUT(n16549), .S0(n102_adj_5275), .S1(n99_adj_5274));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_28 (.A0(d4[61]), .B0(d3[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[62]), .B1(d3[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16547), .COUT(n16548), .S0(n108_adj_5277), .S1(n105_adj_5276));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_28.INJECT1_1 = "NO";
    CCU2C add_4107_17 (.A0(phase_inc_carrGen[14]), .B0(n13099), .C0(n2378), 
          .D0(n18136), .A1(phase_inc_carrGen[15]), .B1(n13099), .C1(n2377), 
          .D1(n3720), .CIN(n16726), .COUT(n16727), .S0(n281), .S1(n278));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_17.INIT0 = 16'h74b8;
    defparam add_4107_17.INIT1 = 16'h74b8;
    defparam add_4107_17.INJECT1_0 = "NO";
    defparam add_4107_17.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_16 (.A0(d_d9_adj_5685[49]), .B0(d9_adj_5684[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[50]), .B1(d9_adj_5684[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16501), .COUT(n16502));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_26 (.A0(d4[59]), .B0(d3[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[60]), .B1(d3[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16546), .COUT(n16547), .S0(n114_adj_5279), .S1(n111_adj_5278));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_24 (.A0(d4[57]), .B0(d3[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[58]), .B1(d3[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16545), .COUT(n16546), .S0(n120_adj_5281), .S1(n117_adj_5280));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_24.INJECT1_1 = "NO";
    CCU2C add_4107_15 (.A0(phase_inc_carrGen[12]), .B0(n13099), .C0(n2380), 
          .D0(n18136), .A1(phase_inc_carrGen[13]), .B1(n13099), .C1(n2379), 
          .D1(n3716), .CIN(n16725), .COUT(n16726), .S0(n287), .S1(n284));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_15.INIT0 = 16'h74b8;
    defparam add_4107_15.INIT1 = 16'h74b8;
    defparam add_4107_15.INJECT1_0 = "NO";
    defparam add_4107_15.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_22 (.A0(d4[55]), .B0(d3[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[56]), .B1(d3[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16544), .COUT(n16545), .S0(n126_adj_5283), .S1(n123_adj_5282));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_20 (.A0(d4[53]), .B0(d3[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[54]), .B1(d3[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16543), .COUT(n16544), .S0(n132_adj_5285), .S1(n129_adj_5284));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_20.INJECT1_1 = "NO";
    CCU2C add_4107_13 (.A0(phase_inc_carrGen[10]), .B0(n13099), .C0(n2382), 
          .D0(n3716), .A1(phase_inc_carrGen[11]), .B1(n13099), .C1(n12207), 
          .D1(n3715), .CIN(n16724), .COUT(n16725), .S0(n293), .S1(n290));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_13.INIT0 = 16'h74b8;
    defparam add_4107_13.INIT1 = 16'h74b8;
    defparam add_4107_13.INJECT1_0 = "NO";
    defparam add_4107_13.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_18 (.A0(d4[51]), .B0(d3[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[52]), .B1(d3[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16542), .COUT(n16543), .S0(n138_adj_5287), .S1(n135_adj_5286));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_16 (.A0(d4[49]), .B0(d3[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[50]), .B1(d3[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16541), .COUT(n16542), .S0(n144_adj_5289), .S1(n141_adj_5288));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_16.INJECT1_1 = "NO";
    CCU2C add_4107_11 (.A0(phase_inc_carrGen[8]), .B0(n13099), .C0(n2384), 
          .D0(n3685), .A1(phase_inc_carrGen[9]), .B1(n13099), .C1(n2383), 
          .D1(n18131), .CIN(n16723), .COUT(n16724), .S0(n299), .S1(n296));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_11.INIT0 = 16'h74b8;
    defparam add_4107_11.INIT1 = 16'h74b8;
    defparam add_4107_11.INJECT1_0 = "NO";
    defparam add_4107_11.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_14 (.A0(d4[47]), .B0(d3[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[48]), .B1(d3[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16540), .COUT(n16541), .S0(n150_adj_5291), .S1(n147_adj_5290));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_12 (.A0(d4[45]), .B0(d3[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[46]), .B1(d3[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16539), .COUT(n16540), .S0(n156_adj_5293), .S1(n153_adj_5292));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_12.INJECT1_1 = "NO";
    CCU2C add_4107_9 (.A0(phase_inc_carrGen[6]), .B0(n13099), .C0(n2386), 
          .D0(n3720), .A1(phase_inc_carrGen[7]), .B1(n13099), .C1(n2385), 
          .D1(n18131), .CIN(n16722), .COUT(n16723), .S0(n305), .S1(n302));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_9.INIT0 = 16'h74b8;
    defparam add_4107_9.INIT1 = 16'h74b8;
    defparam add_4107_9.INJECT1_0 = "NO";
    defparam add_4107_9.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_10 (.A0(d4[43]), .B0(d3[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[44]), .B1(d3[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16538), .COUT(n16539), .S0(n162_adj_5295), .S1(n159_adj_5294));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_8 (.A0(d4[41]), .B0(d3[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[42]), .B1(d3[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16537), .COUT(n16538), .S0(n168_adj_5297), .S1(n165_adj_5296));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_6 (.A0(d4[39]), .B0(d3[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[40]), .B1(d3[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16536), .COUT(n16537), .S0(n174_adj_5299), .S1(n171_adj_5298));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_6.INJECT1_1 = "NO";
    CCU2C add_4107_7 (.A0(phase_inc_carrGen[4]), .B0(n13099), .C0(n2388), 
          .D0(n3720), .A1(phase_inc_carrGen[5]), .B1(n13099), .C1(n2387), 
          .D1(n3720), .CIN(n16721), .COUT(n16722), .S0(n311), .S1(n308));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(256[2] 283[5])
    defparam add_4107_7.INIT0 = 16'h74b8;
    defparam add_4107_7.INIT1 = 16'h74b8;
    defparam add_4107_7.INJECT1_0 = "NO";
    defparam add_4107_7.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_36 (.A0(d_d9_adj_5685[69]), .B0(d9_adj_5684[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5685[70]), .B1(d9_adj_5684[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16511), .COUT(n16512), .S0(n84_adj_4911), 
          .S1(n81_adj_4910));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam _add_1_1637_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_4 (.A0(d4[37]), .B0(d3[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[38]), .B1(d3[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16535), .COUT(n16536), .S0(n180_adj_5301), .S1(n177_adj_5300));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(68[13:20])
    defparam _add_1_1562_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_4.INJECT1_1 = "NO";
    \CIC(width=72,decimation_ratio=4096)_U1  CIC1Cos (.d_d8({d_d8_adj_5683}), 
            .n3(n3_adj_4615), .d_tmp({d_tmp_adj_5671}), .clk_80mhz(clk_80mhz), 
            .d5({d5_adj_5677}), .d_d_tmp({d_d_tmp_adj_5672}), .d2({d2_adj_5674}), 
            .d2_71__N_490({d2_71__N_490_adj_5690}), .d3({d3_adj_5675}), 
            .d3_71__N_562({d3_71__N_562_adj_5691}), .d4({d4_adj_5676}), 
            .d4_71__N_634({d4_71__N_634_adj_5692}), .d5_71__N_706({d5_71__N_706_adj_5693}), 
            .d6({d6_adj_5678}), .d6_71__N_1459({d6_71__N_1459_adj_5705}), 
            .d_d6({d_d6_adj_5679}), .d7({d7_adj_5680}), .d7_71__N_1531({d7_71__N_1531_adj_5706}), 
            .d_d7({d_d7_adj_5681}), .d8({d8_adj_5682}), .d8_71__N_1603({d8_71__N_1603_adj_5707}), 
            .d9({d9_adj_5684}), .d9_71__N_1675({d9_71__N_1675_adj_5708}), 
            .d_d9({d_d9_adj_5685}), .CIC1_outCos({CIC1_outCos}), .d1({d1_adj_5673}), 
            .d1_71__N_418({d1_71__N_418_adj_5689}), .n15(n15_adj_4679), 
            .count({count_adj_5688}), .n28(n28_adj_2750), .n14(n14_adj_4680), 
            .n2(n2_adj_4616), .n87_adj_114({n36_adj_5151, n39_adj_5152, 
            n42_adj_5153, n45_adj_5154, n48_adj_5155, n51_adj_5156, 
            n54_adj_5157, n57_adj_5158, n60_adj_5159, n63_adj_5160, 
            n66_adj_5161, n69_adj_5162, n72_adj_5163, n75_adj_5164, 
            n78_adj_5165, n81_adj_5166}), .n17(n17_adj_4677), .n3_adj_1(n3_adj_4653), 
            .n9(n9), .n2_adj_2(n2_adj_4654), .n5(n5_adj_4651), .n8(n8), 
            .n4(n4_adj_4652), .n7(n7_adj_4649), .n23(n23_adj_4595), .n22(n22_adj_4596), 
            .n2_adj_3(n2_adj_2761), .n25(n25_adj_4593), .n5_adj_4(n5_adj_2758), 
            .n4_adj_5(n4_adj_2759), .\CICGain[1] (CICGain[1]), .\d10[60] (d10_adj_5686[60]), 
            .n17784(n17784), .\d10[59] (d10_adj_5686[59]), .n24(n24_adj_4594), 
            .n27(n27_adj_4588), .n26(n26_adj_4589), .n29(n29_adj_4586), 
            .n28_adj_6(n28_adj_4587), .n31(n31_adj_4584), .n30(n30_adj_4585), 
            .n7_adj_7(n7_adj_2756), .n33(n33_adj_4582), .n6(n6_adj_4650), 
            .n6_adj_8(n6_adj_2757), .n11(n11), .n10(n10), .n32(n32_adj_4583), 
            .n9_adj_9(n9_adj_4647), .n8_adj_10(n8_adj_4648), .n35(n35_adj_4580), 
            .n34(n34_adj_4581), .n17805(n17805), .\d10[62] (d10_adj_5686[62]), 
            .\d10[63] (d10_adj_5686[63]), .\CICGain[0] (CICGain[0]), .n63_adj_11(n63), 
            .n37(n37_adj_4578), .n29_adj_12(n29_adj_2749), .n5_adj_13(n5_adj_4613), 
            .n36_adj_14(n36_adj_4579), .n16(n16_adj_4678), .n13(n13), 
            .n12(n12), .n15_adj_15(n15), .n14_adj_16(n14), .n17_adj_17(n17), 
            .n16_adj_18(n16), .n19(n19), .n18(n18), .n21(n21), .n20(n20), 
            .\d10[61] (d10_adj_5686[61]), .\d10[64] (d10_adj_5686[64]), 
            .\d10[65] (d10_adj_5686[65]), .\d10[66] (d10_adj_5686[66]), 
            .\d10[67] (d10_adj_5686[67]), .\d10[68] (d10_adj_5686[68]), 
            .\d10[69] (d10_adj_5686[69]), .\d10[70] (d10_adj_5686[70]), 
            .\d10[71] (d10_adj_5686[71]), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_5711[2]), 
            .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_5711[3]), .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_5711[4]), 
            .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_5711[5]), .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_5711[6]), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_5711[7]), .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_5711[8]), 
            .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_5711[9]), .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5711[10]), 
            .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5711[11]), .n19_adj_19(n19_adj_4675), 
            .n11_adj_20(n11_adj_4645), .n33_adj_21(n33), .n32_adj_22(n32), 
            .n35_adj_23(n35), .n10_adj_24(n10_adj_4646), .n13_adj_25(n13_adj_4643), 
            .n12_adj_26(n12_adj_4644), .n15_adj_27(n15_adj_4641), .n14_adj_28(n14_adj_4642), 
            .n17_adj_29(n17_adj_4639), .n16_adj_30(n16_adj_4640), .n19_adj_31(n19_adj_4637), 
            .n18_adj_32(n18_adj_4638), .n21_adj_33(n21_adj_4635), .n20_adj_34(n20_adj_4636), 
            .n23_adj_35(n23_adj_4633), .n22_adj_36(n22_adj_4634), .n25_adj_37(n25_adj_4631), 
            .n24_adj_38(n24_adj_4632), .n3_adj_39(n3), .n27_adj_40(n27_adj_4629), 
            .n26_adj_41(n26_adj_4630), .n2_adj_42(n2), .n5_adj_43(n5), 
            .n29_adj_44(n29_adj_4627), .n28_adj_45(n28_adj_4628), .n4_adj_46(n4), 
            .n7_adj_47(n7), .n31_adj_48(n31_adj_4624), .n30_adj_49(n30_adj_4626), 
            .n6_adj_50(n6), .n9_adj_51(n9_adj_4682), .n33_adj_52(n33_adj_4622), 
            .n32_adj_53(n32_adj_4623), .n8_adj_54(n8_adj_4686), .n11_adj_55(n11_adj_4684), 
            .n35_adj_56(n35_adj_4620), .n34_adj_57(n34_adj_4621), .n4_adj_58(n4_adj_4614), 
            .n10_adj_59(n10_adj_4683), .n13_adj_60(n13_adj_4681), .n34_adj_61(n34), 
            .n23_adj_62(n23_adj_2755), .n22_adj_63(n22), .n27_adj_64(n27_adj_2751), 
            .n26_adj_65(n26_adj_2752), .n37_adj_66(n37_adj_4618), .n36_adj_67(n36_adj_4619), 
            .n12_adj_68(n12_adj_4685), .n18_adj_69(n18_adj_4676), .n21_adj_70(n21_adj_4673), 
            .n64(n64), .n7_adj_71(n7_adj_4611), .n65(n65), .n20_adj_72(n20_adj_4674), 
            .n18_adj_73(n18_adj_4600), .n23_adj_74(n23_adj_4671), .n22_adj_75(n22_adj_4672), 
            .n21_adj_76(n21_adj_4597), .n6_adj_77(n6_adj_4612), .n25_adj_78(n25_adj_4669), 
            .n24_adj_79(n24_adj_4670), .n66_adj_80(n66), .n9_adj_81(n9_adj_4609), 
            .n8_adj_82(n8_adj_4610), .n27_adj_83(n27_adj_4667), .n11_adj_84(n11_adj_4607), 
            .n10_adj_85(n10_adj_4608), .n26_adj_86(n26_adj_4668), .n29_adj_87(n29_adj_4665), 
            .n28_adj_88(n28_adj_4666), .n31_adj_89(n31_adj_4663), .n30_adj_90(n30_adj_4664), 
            .n13_adj_91(n13_adj_4605), .n33_adj_92(n33_adj_4661), .n32_adj_93(n32_adj_4662), 
            .n12_adj_94(n12_adj_4606), .n35_adj_95(n35_adj_4659), .n15_adj_96(n15_adj_4603), 
            .n34_adj_97(n34_adj_4660), .n31_adj_98(n31), .n30_adj_99(n30_adj_2748), 
            .n37_adj_100(n37_adj_4656), .n14_adj_101(n14_adj_4604), .n36_adj_102(n36_adj_4657), 
            .n20_adj_103(n20_adj_4598), .n17_adj_104(n17_adj_4601), .n16_adj_105(n16_adj_4602), 
            .n19_adj_106(n19_adj_4599), .n118(n118_adj_5559), .n120(n120_adj_4923), 
            .cout(cout_adj_5229), .n115(n115_adj_5558), .n117(n117_adj_4922), 
            .n112(n112_adj_5557), .n114(n114_adj_4921), .n109(n109_adj_5556), 
            .n111(n111_adj_4920), .n106(n106_adj_5555), .n108(n108_adj_4919), 
            .n37_adj_107(n37), .n36_adj_108(n36), .n103(n103_adj_5554), 
            .n105(n105_adj_4918), .n100(n100_adj_5553), .n102(n102_adj_4917), 
            .n97(n97_adj_5552), .n99(n99_adj_4916), .n94(n94_adj_5551), 
            .n96(n96_adj_4915), .n91(n91_adj_5550), .n93(n93_adj_4914), 
            .n25_adj_109(n25_adj_2753), .n88(n88_adj_5549), .n90(n90_adj_4913), 
            .n24_adj_110(n24_adj_2754), .n85(n85_adj_5548), .n87(n87_adj_4912), 
            .n82(n82_adj_5547), .n84(n84_adj_4911), .n79(n79_adj_5546), 
            .n81_adj_111(n81_adj_4910), .n76(n76_adj_5545), .n78_adj_112(n78_adj_4909), 
            .n3_adj_113(n3_adj_2760)) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(190[45] 196[2])
    AMDemodulator AMDemodulator1 (.\d_out_d_11__N_1892[17] (d_out_d_11__N_1892[17]), 
            .CIC1_out_clkSin(CIC1_out_clkSin), .CIC1_outSin({CIC1_outSin}), 
            .CIC1_outCos({CIC1_outCos}), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
            .\d_out_d_11__N_1890[17] (d_out_d_11__N_1890[17]), .\d_out_d_11__N_1888[17] (d_out_d_11__N_1888[17]), 
            .\d_out_d_11__N_1886[17] (d_out_d_11__N_1886[17]), .\d_out_d_11__N_1884[17] (d_out_d_11__N_1884[17]), 
            .\d_out_d_11__N_1882[17] (d_out_d_11__N_1882[17]), .\d_out_d_11__N_1880[17] (d_out_d_11__N_1880[17]), 
            .d_out_d_11__N_1879(d_out_d_11__N_1879), .\d_out_d_11__N_1878[17] (d_out_d_11__N_1878[17]), 
            .d_out_d_11__N_1877(d_out_d_11__N_1877), .\d_out_d_11__N_1876[17] (d_out_d_11__N_1876[17]), 
            .d_out_d_11__N_1875(d_out_d_11__N_1875), .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), 
            .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), 
            .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), 
            .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), 
            .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DemodOut[9] (DemodOut[9]), 
            .\ISquare[31] (ISquare[31]), .n209(n209), .\d_out_d_11__N_2335[17] (d_out_d_11__N_2335[17]), 
            .\d_out_d_11__N_2353[17] (d_out_d_11__N_2353[17]), .\d_out_d_11__N_1874[17] (d_out_d_11__N_1874[17]), 
            .d_out_d_11__N_1873(d_out_d_11__N_1873), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultResult2({MultResult2}), .MultResult1({MultResult1})) /* synthesis syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(222[15] 227[10])
    LUT4 i1_2_lut_rep_168_3_lut_4_lut (.A(led_c_1), .B(led_c_4), .C(n26_adj_5659), 
         .D(led_c_0), .Z(n18138)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_168_3_lut_4_lut.init = 16'h0020;
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (MixerOutSin, clk_80mhz, DiffOut_c, MixerOutCos, RFIn_c, 
            \LOSine[2] , MixerOutSin_11__N_236, \LOSine[3] , \LOSine[4] , 
            \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , \LOSine[9] , 
            \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[2] , 
            MixerOutCos_11__N_250, \LOCosine[3] , \LOCosine[1] , \LOCosine[4] , 
            \LOCosine[5] , \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , 
            \LOCosine[9] , \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , 
            \LOSine[1] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]MixerOutSin;
    input clk_80mhz;
    output DiffOut_c;
    output [11:0]MixerOutCos;
    input RFIn_c;
    input \LOSine[2] ;
    input [11:0]MixerOutSin_11__N_236;
    input \LOSine[3] ;
    input \LOSine[4] ;
    input \LOSine[5] ;
    input \LOSine[6] ;
    input \LOSine[7] ;
    input \LOSine[8] ;
    input \LOSine[9] ;
    input \LOSine[10] ;
    input \LOSine[11] ;
    input \LOSine[12] ;
    input \LOCosine[2] ;
    input [11:0]MixerOutCos_11__N_250;
    input \LOCosine[3] ;
    input \LOCosine[1] ;
    input \LOCosine[4] ;
    input \LOCosine[5] ;
    input \LOCosine[6] ;
    input \LOCosine[7] ;
    input \LOCosine[8] ;
    input \LOCosine[9] ;
    input \LOCosine[10] ;
    input \LOCosine[11] ;
    input \LOCosine[12] ;
    input \LOSine[1] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    wire [11:0]MixerOutSin_11__N_212;
    
    wire RFInR;
    wire [11:0]MixerOutCos_11__N_224;
    
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_212[0]), .CK(clk_80mhz), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(clk_80mhz), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(23[10] 27[8])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_224[0]), .CK(clk_80mhz), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(clk_80mhz), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(23[10] 27[8])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_212[1]), .CK(clk_80mhz), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_212[2]), .CK(clk_80mhz), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_212[3]), .CK(clk_80mhz), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_212[4]), .CK(clk_80mhz), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_212[5]), .CK(clk_80mhz), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_212[6]), .CK(clk_80mhz), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_212[7]), .CK(clk_80mhz), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_212[8]), .CK(clk_80mhz), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_212[9]), .CK(clk_80mhz), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_212[10]), .CK(clk_80mhz), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_212[11]), .CK(clk_80mhz), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_224[1]), .CK(clk_80mhz), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_224[2]), .CK(clk_80mhz), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_224[3]), .CK(clk_80mhz), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_224[4]), .CK(clk_80mhz), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_224[5]), .CK(clk_80mhz), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_224[6]), .CK(clk_80mhz), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_224[7]), .CK(clk_80mhz), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_224[8]), .CK(clk_80mhz), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_224[9]), .CK(clk_80mhz), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_224[10]), .CK(clk_80mhz), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_224[11]), .CK(clk_80mhz), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=170, LSE_RLINE=178 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_236[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_236[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_236[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_236[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_236[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_236[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_236[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_236[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_236[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_236[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_236[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_250[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_250[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_250[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_250[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_250[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_250[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_250[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_250[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_250[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_250[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_250[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_250[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_236[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (\DemodOut[9] , \DataInReg[0] , clk_80mhz, \DataInReg_11__N_1856[0] , 
            counter, GND_net, VCC_net, \DataInReg[1] , \DataInReg_11__N_1856[1] , 
            \DataInReg[2] , \DataInReg_11__N_1856[2] , \DataInReg[3] , 
            \DataInReg_11__N_1856[3] , \DataInReg[4] , \DataInReg_11__N_1856[4] , 
            \DataInReg[5] , \DataInReg_11__N_1856[5] , \DataInReg[6] , 
            \DataInReg_11__N_1856[6] , \DataInReg[7] , \DataInReg_11__N_1856[7] , 
            \DataInReg[8] , \DataInReg_11__N_1856[8] , \DataInReg[9] ) /* synthesis syn_module_defined=1 */ ;
    input \DemodOut[9] ;
    output \DataInReg[0] ;
    input clk_80mhz;
    input \DataInReg_11__N_1856[0] ;
    output [9:0]counter;
    input GND_net;
    input VCC_net;
    output \DataInReg[1] ;
    input \DataInReg_11__N_1856[1] ;
    output \DataInReg[2] ;
    input \DataInReg_11__N_1856[2] ;
    output \DataInReg[3] ;
    input \DataInReg_11__N_1856[3] ;
    output \DataInReg[4] ;
    input \DataInReg_11__N_1856[4] ;
    output \DataInReg[5] ;
    input \DataInReg_11__N_1856[5] ;
    output \DataInReg[6] ;
    input \DataInReg_11__N_1856[6] ;
    output \DataInReg[7] ;
    input \DataInReg_11__N_1856[7] ;
    output \DataInReg[8] ;
    input \DataInReg_11__N_1856[8] ;
    output \DataInReg[9] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    wire [11:0]n3976;
    
    wire clk_80mhz_enable_1469, n16715;
    wire [9:0]n45;
    
    wire n16714, n16713, n16712, n16711, n17, n15, n11, n12;
    
    LUT4 i1156_1_lut (.A(\DemodOut[9] ), .Z(n3976[9])) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(26[3] 27[35])
    defparam i1156_1_lut.init = 16'h5555;
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1856[0] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i1.GSR = "ENABLED";
    CCU2C counter_1006_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16715), .S0(n45[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_11.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_11.INIT1 = 16'h0000;
    defparam counter_1006_add_4_11.INJECT1_0 = "NO";
    defparam counter_1006_add_4_11.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16714), .COUT(n16715), .S0(n45[7]), .S1(n45[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_9.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_9.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_9.INJECT1_0 = "NO";
    defparam counter_1006_add_4_9.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16713), .COUT(n16714), .S0(n45[5]), .S1(n45[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_7.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_7.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_7.INJECT1_0 = "NO";
    defparam counter_1006_add_4_7.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16712), .COUT(n16713), .S0(n45[3]), .S1(n45[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_5.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_5.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_5.INJECT1_0 = "NO";
    defparam counter_1006_add_4_5.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16711), .COUT(n16712), .S0(n45[1]), .S1(n45[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_3.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_3.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_3.INJECT1_0 = "NO";
    defparam counter_1006_add_4_3.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16711), .S1(n45[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_1.INIT0 = 16'h0000;
    defparam counter_1006_add_4_1.INIT1 = 16'h555f;
    defparam counter_1006_add_4_1.INJECT1_0 = "NO";
    defparam counter_1006_add_4_1.INJECT1_1 = "NO";
    FD1S3AX counter_1006__i0 (.D(n45[0]), .CK(clk_80mhz), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i0.GSR = "ENABLED";
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1856[1] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1856[2] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1856[3] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1856[4] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1856[5] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1856[6] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1856[7] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1856[8] ), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(\DataInReg[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n3976[9]), .SP(clk_80mhz_enable_1469), .CK(clk_80mhz), 
            .Q(\DataInReg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=199, LSE_RLINE=205 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i10.GSR = "ENABLED";
    LUT4 i6638_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(clk_80mhz_enable_1469)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(26[7:19])
    defparam i6638_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(26[7:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(counter[6]), .B(counter[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(26[7:19])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(26[7:19])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[8]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(26[7:19])
    defparam i2_2_lut.init = 16'heeee;
    FD1S3AX counter_1006__i1 (.D(n45[1]), .CK(clk_80mhz), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i1.GSR = "ENABLED";
    FD1S3AX counter_1006__i2 (.D(n45[2]), .CK(clk_80mhz), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i2.GSR = "ENABLED";
    FD1S3AX counter_1006__i3 (.D(n45[3]), .CK(clk_80mhz), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i3.GSR = "ENABLED";
    FD1S3AX counter_1006__i4 (.D(n45[4]), .CK(clk_80mhz), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i4.GSR = "ENABLED";
    FD1S3AX counter_1006__i5 (.D(n45[5]), .CK(clk_80mhz), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i5.GSR = "ENABLED";
    FD1S3AX counter_1006__i6 (.D(n45[6]), .CK(clk_80mhz), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i6.GSR = "ENABLED";
    FD1S3AX counter_1006__i7 (.D(n45[7]), .CK(clk_80mhz), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i7.GSR = "ENABLED";
    FD1S3AX counter_1006__i8 (.D(n45[8]), .CK(clk_80mhz), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i8.GSR = "ENABLED";
    FD1S3AX counter_1006__i9 (.D(n45[9]), .CK(clk_80mhz), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/PWM.v(25[14:29])
    defparam counter_1006__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (clk_80mhz, i_Rx_Serial_c, o_Rx_Byte1, 
            GND_net, VCC_net, o_Rx_DV1) /* synthesis syn_module_defined=1 */ ;
    input clk_80mhz;
    input i_Rx_Serial_c;
    output [7:0]o_Rx_Byte1;
    input GND_net;
    input VCC_net;
    output o_Rx_DV1;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx1/UartClk[2], is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(37[14:21])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    wire [2:0]r_SM_Main;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(43[17:26])
    wire [2:0]r_SM_Main_2__N_2424;
    
    wire n17609, UartClk_2_enable_30, n18034, r_Rx_DV_last, r_Rx_DV, 
        r_Rx_Data_R, r_Rx_Data, UartClk_2_enable_15;
    wire [7:0]r_Rx_Byte;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(41[17:26])
    
    wire UartClk_2_enable_2, n16709;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire n16708;
    wire [15:0]r_Clock_Count;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(39[18:31])
    wire [15:0]n69;
    wire [2:0]r_Bit_Index;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(40[17:28])
    
    wire UartClk_2_enable_32, n17446, n17394, n18140, n12631, n16707, 
        n16706, n18133, n17326, n17269, n13103, n18163, n18162, 
        UartClk_2_enable_5, n18148, n18128, n16705, n12996, n18032, 
        r_Rx_DV_N_2484, n18130, n17313, UartClk_2_enable_6, n16704, 
        n16703, UartClk_2_enable_4, n17300, UartClk_2_enable_7;
    wire [2:0]n132;
    
    wire n17449, n16702, n16701, n18164, n17740, n17601, n26, 
        n17491, n17587, UartClk_2_enable_35, UartClk_2_enable_34, n18033, 
        n12615, r_Rx_DV_last_N_2483, UartClk_2_enable_36, UartClk_2_enable_33, 
        n13079, n17579, n17581, n17573, n17577;
    
    LUT4 i6630_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main_2__N_2424[0]), 
         .D(n17609), .Z(UartClk_2_enable_30)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i6630_4_lut.init = 16'h5455;
    FD1S3IX r_SM_Main_i0 (.D(n18034), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(clk_80mhz), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_2), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    CCU2C UartClk_1007_1031_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16709), .S0(n17[1]), .S1(n17[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031_add_4_3.INIT0 = 16'haaa0;
    defparam UartClk_1007_1031_add_4_3.INIT1 = 16'haaa0;
    defparam UartClk_1007_1031_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_1007_1031_add_4_3.INJECT1_1 = "NO";
    CCU2C UartClk_1007_1031_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16709), .S1(n17[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031_add_4_1.INIT0 = 16'h0000;
    defparam UartClk_1007_1031_add_4_1.INIT1 = 16'h555f;
    defparam UartClk_1007_1031_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_1007_1031_add_4_1.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16708), .S0(n69[15]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_17.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_1009_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_17.INJECT1_1 = "NO";
    FD1P3AX r_Bit_Index_i0 (.D(n17446), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n17609)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(r_SM_Main[2]), .B(n17394), .C(n18140), .D(r_SM_Main[1]), 
         .Z(n12631)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h5011;
    LUT4 i6184_3_lut (.A(r_SM_Main[0]), .B(r_Rx_Data), .C(r_SM_Main_2__N_2424[0]), 
         .Z(n17394)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i6184_3_lut.init = 16'ha8a8;
    CCU2C r_Clock_Count_1009_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16707), .COUT(n16708), .S0(n69[13]), 
          .S1(n69[14]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_15.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_15.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_15.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16706), .COUT(n16707), .S0(n69[11]), 
          .S1(n69[12]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_13.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_13.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_13.INJECT1_1 = "NO";
    LUT4 i6607_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n18133), .C(n17326), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_2)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i6607_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(r_SM_Main[0]), 
         .B(n17269), .C(n13103), .Z(n18163)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h5757;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main[0]), 
         .B(r_SM_Main_2__N_2424[0]), .C(r_Rx_Data), .Z(n18162)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_rep_170 (.A(n13103), .B(n17269), .Z(n18140)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_170.init = 16'heeee;
    LUT4 i6601_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n18133), .C(n17326), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_5)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i6601_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i6632_2_lut_3_lut_4_lut (.A(n13103), .B(n17269), .C(r_SM_Main[0]), 
         .D(n18148), .Z(UartClk_2_enable_15)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i6632_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_rep_158_3_lut_4_lut (.A(n13103), .B(n17269), .C(r_SM_Main[0]), 
         .D(n18148), .Z(n18128)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_158_3_lut_4_lut.init = 16'hfff1;
    CCU2C r_Clock_Count_1009_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16705), .COUT(n16706), .S0(n69[9]), 
          .S1(n69[10]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_11.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_11.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_11.INJECT1_1 = "NO";
    LUT4 r_SM_Main_2__N_2418_2__bdd_3_lut_6652_4_lut (.A(n13103), .B(n17269), 
         .C(r_SM_Main[0]), .D(n12996), .Z(n18032)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam r_SM_Main_2__N_2418_2__bdd_3_lut_6652_4_lut.init = 16'h1e10;
    LUT4 i6589_2_lut_3_lut_4_lut (.A(n13103), .B(n17269), .C(n18148), 
         .D(r_SM_Main[0]), .Z(r_Rx_DV_N_2484)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i6589_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i2351_2_lut_rep_160_3_lut (.A(n13103), .B(n17269), .C(r_SM_Main[0]), 
         .Z(n18130)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i2351_2_lut_rep_160_3_lut.init = 16'hf1f1;
    LUT4 i6578_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n18133), .C(n17313), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_6)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i6578_2_lut_3_lut_4_lut.init = 16'h0001;
    CCU2C r_Clock_Count_1009_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16704), .COUT(n16705), .S0(n69[7]), 
          .S1(n69[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_9.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_9.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_9.INJECT1_1 = "NO";
    FD1S3AX UartClk_1007_1031__i0 (.D(n17[0]), .CK(clk_80mhz), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031__i0.GSR = "ENABLED";
    CCU2C r_Clock_Count_1009_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16703), .COUT(n16704), .S0(n69[5]), 
          .S1(n69[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_7.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_7.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_7.INJECT1_1 = "NO";
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_4), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_5), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_6), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(n18140), .CK(UartClk[2]), .CD(n17300), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2484), .SP(UartClk_2_enable_7), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_45 (.A(n132[2]), .B(n18130), .C(n12996), .D(r_SM_Main[1]), 
         .Z(n17449)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_45.init = 16'h0200;
    CCU2C r_Clock_Count_1009_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16702), .COUT(n16703), .S0(n69[3]), 
          .S1(n69[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_5.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_5.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_5.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16701), .COUT(n16702), .S0(n69[1]), 
          .S1(n69[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_3.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_3.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_3.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16701), .S1(n69[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_1.INIT0 = 16'h0000;
    defparam r_Clock_Count_1009_add_4_1.INIT1 = 16'h555f;
    defparam r_Clock_Count_1009_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_1.INJECT1_1 = "NO";
    FD1S3IX r_SM_Main_i1 (.D(n18164), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i0 (.D(n69[0]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i0.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[4]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[6]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i1173_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), .C(r_Bit_Index[0]), 
         .Z(n132[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(119[36:54])
    defparam i1173_3_lut.init = 16'h6a6a;
    LUT4 i1_4_lut_adj_46 (.A(n17740), .B(n17269), .C(n17601), .D(r_Clock_Count[1]), 
         .Z(r_SM_Main_2__N_2424[0])) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i1_4_lut_adj_46.init = 16'hfdff;
    LUT4 i6528_2_lut (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), .Z(n17740)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6528_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_47 (.A(n26), .B(n18140), .C(r_SM_Main[0]), .D(r_SM_Main[1]), 
         .Z(n17491)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_47.init = 16'h0800;
    LUT4 i39_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n26)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i39_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_48 (.A(r_Clock_Count[0]), .B(r_Clock_Count[6]), .C(r_Clock_Count[2]), 
         .D(r_Clock_Count[4]), .Z(n17601)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_48.init = 16'hfffd;
    LUT4 i1_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[0]), .C(r_Bit_Index[1]), 
         .Z(n12996)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i6575_4_lut (.A(n17587), .B(n17269), .C(n13103), .D(r_SM_Main[1]), 
         .Z(UartClk_2_enable_32)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i6575_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_49 (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .Z(n17587)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_49.init = 16'heeee;
    LUT4 i6612_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n18128), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_35)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(114[17:39])
    defparam i6612_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i6615_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n18128), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_34)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(114[17:39])
    defparam i6615_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 r_SM_Main_2__N_2418_2__bdd_3_lut (.A(r_SM_Main_2__N_2424[0]), .B(r_Rx_Data), 
         .C(r_SM_Main[0]), .Z(n18033)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(C))) */ ;
    defparam r_SM_Main_2__N_2418_2__bdd_3_lut.init = 16'ha3a3;
    LUT4 i1_2_lut_adj_50 (.A(r_Bit_Index[0]), .B(r_Bit_Index[2]), .Z(n17313)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(114[17:39])
    defparam i1_2_lut_adj_50.init = 16'heeee;
    FD1P3IX r_Clock_Count_1009__i15 (.D(n69[15]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i15.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_178 (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .Z(n18148)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_178.init = 16'hbbbb;
    LUT4 i2878_1_lut (.A(r_Rx_DV), .Z(n12615)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i2878_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2483)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_163_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), 
         .C(n17269), .D(n13103), .Z(n18133)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i1_2_lut_rep_163_3_lut_4_lut.init = 16'hbbbf;
    LUT4 i6610_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n18128), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(114[17:39])
    defparam i6610_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i6617_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n18128), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_33)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(114[17:39])
    defparam i6617_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i6598_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n17300)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i6598_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(n18140), .Z(UartClk_2_enable_7)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i21_4_lut_4_lut.init = 16'h2505;
    LUT4 i3366_4_lut (.A(n13079), .B(r_Clock_Count[6]), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[4]), .Z(n13103)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i3366_4_lut.init = 16'hc8c0;
    LUT4 i3342_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n13079)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i3342_3_lut.init = 16'hecec;
    PFUMX i6653 (.BLUT(n18033), .ALUT(n18032), .C0(r_SM_Main[1]), .Z(n18034));
    LUT4 i1_4_lut_adj_51 (.A(n17579), .B(n17581), .C(n17573), .D(n17577), 
         .Z(n17269)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_51.init = 16'hfffe;
    FD1S3AX UartClk_1007_1031__i1 (.D(n17[1]), .CK(clk_80mhz), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031__i1.GSR = "ENABLED";
    FD1S3AX UartClk_1007_1031__i2 (.D(n17[2]), .CK(clk_80mhz), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031__i2.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_52 (.A(r_Clock_Count[11]), .B(r_Clock_Count[15]), 
         .Z(n17579)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_52.init = 16'heeee;
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2483), .CK(clk_80mhz), .CD(n12615), 
            .Q(o_Rx_DV1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i14 (.D(n69[14]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i14.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i13 (.D(n69[13]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i13.GSR = "ENABLED";
    LUT4 i1_3_lut_adj_53 (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), .C(r_Clock_Count[7]), 
         .Z(n17581)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_3_lut_adj_53.init = 16'hfefe;
    FD1P3IX r_Clock_Count_1009__i12 (.D(n69[12]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i12.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_54 (.A(r_Clock_Count[14]), .B(r_Clock_Count[10]), 
         .Z(n17573)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_54.init = 16'heeee;
    FD1P3IX r_Clock_Count_1009__i11 (.D(n69[11]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i11.GSR = "ENABLED";
    LUT4 i6645_3_lut_4_lut (.A(n18140), .B(r_SM_Main[0]), .C(r_Bit_Index[0]), 
         .D(r_SM_Main[1]), .Z(n17446)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i6645_3_lut_4_lut.init = 16'h0200;
    LUT4 i6604_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n18133), .C(n17313), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_4)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i6604_2_lut_3_lut_4_lut.init = 16'h0100;
    FD1P3IX r_Clock_Count_1009__i10 (.D(n69[10]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i9 (.D(n69[9]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i9.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_55 (.A(r_Clock_Count[9]), .B(r_Clock_Count[12]), .Z(n17577)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_55.init = 16'heeee;
    FD1P3IX r_Clock_Count_1009__i8 (.D(n69[8]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i7 (.D(n69[7]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i6 (.D(n69[6]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i6.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i5 (.D(n69[5]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i4 (.D(n69[4]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i3 (.D(n69[3]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i2 (.D(n69[2]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i1 (.D(n69[1]), .SP(UartClk_2_enable_30), 
            .CD(n12631), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i1.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i2 (.D(n17449), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n17491), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_56 (.A(r_Bit_Index[2]), .B(r_Bit_Index[0]), .Z(n17326)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(114[17:39])
    defparam i1_2_lut_adj_56.init = 16'hbbbb;
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_33), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_34), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_35), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=230, LSE_RLINE=235 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    PFUMX i6702 (.BLUT(n18162), .ALUT(n18163), .C0(r_SM_Main[1]), .Z(n18164));
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096) 
//

module \CIC(width=72,decimation_ratio=4096)  (d_tmp, clk_80mhz, d5, d_d_tmp, 
            d2, d2_71__N_490, d3, d3_71__N_562, d4, d4_71__N_634, 
            d5_71__N_706, d6, d6_71__N_1459, d_d6, CIC1_out_clkSin, 
            d7, d7_71__N_1531, d_d7, d8, d8_71__N_1603, d_d8, d9, 
            d9_71__N_1675, d_d9, CIC1_outSin, d1, d1_71__N_418, count, 
            n32, n25, n24, \CICGain[1] , \CICGain[0] , n9, n8, 
            n33, n27, n26, n26_adj_115, n32_adj_116, n29, n35, 
            n35_adj_117, \d10[69] , \d10[68] , n34, \d10[65] , \d10[66] , 
            \d10[67] , n11, n10, n37, n36, n28, \d10[70] , \d10[71] , 
            n37_adj_118, n34_adj_119, n37_adj_120, n33_adj_121, n32_adj_122, 
            n36_adj_123, n31, n30, n87_adj_228, n63_adj_125, \d_out_11__N_1819[2] , 
            n5, n11_adj_126, n10_adj_127, n13, n12, n15, n4, n14, 
            n17, n16, n25_adj_128, n24_adj_129, n29_adj_130, n28_adj_131, 
            n31_adj_132, n30_adj_133, n64, \d_out_11__N_1819[3] , n36_adj_134, 
            n65, \d_out_11__N_1819[4] , n66_adj_135, \d_out_11__N_1819[5] , 
            \d_out_11__N_1819[6] , n13_adj_136, n12_adj_137, \d10[64] , 
            n15_adj_138, \d10[62] , \d10[63] , n17784, \d10[60] , 
            n14_adj_139, n17_adj_140, \d10[61] , n17805, \d10[59] , 
            n16_adj_141, n3, n2, n19, n5_adj_142, n4_adj_143, n7, 
            n6, \d_out_11__N_1819[7] , n33_adj_144, n22, n6_adj_145, 
            n19_adj_146, n27_adj_147, n26_adj_148, n29_adj_149, n18, 
            n23, n22_adj_150, n28_adj_151, n21, n20, n18_adj_152, 
            n31_adj_153, n35_adj_154, n34_adj_155, n30_adj_156, n33_adj_157, 
            n25_adj_158, n118, n120, cout, n32_adj_159, n24_adj_160, 
            n115, n117, n35_adj_161, n27_adj_162, n34_adj_163, n26_adj_164, 
            n29_adj_165, n112, n114, n3_adj_166, n109, n111, n106, 
            n108, n103, n105, n37_adj_167, n28_adj_168, n100, n102, 
            n97, n99, n36_adj_169, n94, n96, n91, n93, n88, 
            n90, n2_adj_170, n85, n87, n3_adj_171, n2_adj_172, n5_adj_173, 
            n4_adj_174, n7_adj_175, n82, n84, n6_adj_176, n9_adj_177, 
            n3_adj_178, n8_adj_179, n23_adj_180, n7_adj_181, n2_adj_182, 
            n5_adj_183, n79, n81_adj_184, n9_adj_185, n76, n78_adj_186, 
            n4_adj_187, n11_adj_188, n10_adj_189, n7_adj_190, n6_adj_191, 
            n31_adj_192, n9_adj_193, n21_adj_194, n20_adj_195, n8_adj_196, 
            \d_out_11__N_1819[10] , n11_adj_197, n13_adj_198, n12_adj_199, 
            n30_adj_200, n10_adj_201, n13_adj_202, \d_out_11__N_1819[11] , 
            n8_adj_203, n12_adj_204, n15_adj_205, n15_adj_206, n14_adj_207, 
            n14_adj_208, n17_adj_209, n16_adj_210, n19_adj_211, n17_adj_212, 
            n18_adj_213, n16_adj_214, n21_adj_215, n20_adj_216, n19_adj_217, 
            n23_adj_218, n22_adj_219, n25_adj_220, n18_adj_221, n21_adj_222, 
            n20_adj_223, \d_out_11__N_1819[8] , n24_adj_224, n27_adj_225, 
            n23_adj_226, \d_out_11__N_1819[9] , n22_adj_227) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output CIC1_out_clkSin;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d_d7;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d_d8;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output [11:0]CIC1_outSin;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output [15:0]count;
    output n32;
    output n25;
    output n24;
    input \CICGain[1] ;
    input \CICGain[0] ;
    output n9;
    output n8;
    output n33;
    output n27;
    output n26;
    output n26_adj_115;
    output n32_adj_116;
    output n29;
    output n35;
    output n35_adj_117;
    input \d10[69] ;
    input \d10[68] ;
    output n34;
    input \d10[65] ;
    input \d10[66] ;
    input \d10[67] ;
    output n11;
    output n10;
    output n37;
    output n36;
    output n28;
    input \d10[70] ;
    input \d10[71] ;
    output n37_adj_118;
    output n34_adj_119;
    output n37_adj_120;
    output n33_adj_121;
    output n32_adj_122;
    output n36_adj_123;
    output n31;
    output n30;
    input [15:0]n87_adj_228;
    input n63_adj_125;
    output \d_out_11__N_1819[2] ;
    output n5;
    output n11_adj_126;
    output n10_adj_127;
    output n13;
    output n12;
    output n15;
    output n4;
    output n14;
    output n17;
    output n16;
    output n25_adj_128;
    output n24_adj_129;
    output n29_adj_130;
    output n28_adj_131;
    output n31_adj_132;
    output n30_adj_133;
    input n64;
    output \d_out_11__N_1819[3] ;
    output n36_adj_134;
    input n65;
    output \d_out_11__N_1819[4] ;
    input n66_adj_135;
    output \d_out_11__N_1819[5] ;
    output \d_out_11__N_1819[6] ;
    output n13_adj_136;
    output n12_adj_137;
    input \d10[64] ;
    output n15_adj_138;
    input \d10[62] ;
    input \d10[63] ;
    input n17784;
    input \d10[60] ;
    output n14_adj_139;
    output n17_adj_140;
    input \d10[61] ;
    input n17805;
    input \d10[59] ;
    output n16_adj_141;
    output n3;
    output n2;
    output n19;
    output n5_adj_142;
    output n4_adj_143;
    output n7;
    output n6;
    output \d_out_11__N_1819[7] ;
    output n33_adj_144;
    output n22;
    output n6_adj_145;
    output n19_adj_146;
    output n27_adj_147;
    output n26_adj_148;
    output n29_adj_149;
    output n18;
    output n23;
    output n22_adj_150;
    output n28_adj_151;
    output n21;
    output n20;
    output n18_adj_152;
    output n31_adj_153;
    output n35_adj_154;
    output n34_adj_155;
    output n30_adj_156;
    output n33_adj_157;
    output n25_adj_158;
    input n118;
    input n120;
    input cout;
    output n32_adj_159;
    output n24_adj_160;
    input n115;
    input n117;
    output n35_adj_161;
    output n27_adj_162;
    output n34_adj_163;
    output n26_adj_164;
    output n29_adj_165;
    input n112;
    input n114;
    output n3_adj_166;
    input n109;
    input n111;
    input n106;
    input n108;
    input n103;
    input n105;
    output n37_adj_167;
    output n28_adj_168;
    input n100;
    input n102;
    input n97;
    input n99;
    output n36_adj_169;
    input n94;
    input n96;
    input n91;
    input n93;
    input n88;
    input n90;
    output n2_adj_170;
    input n85;
    input n87;
    output n3_adj_171;
    output n2_adj_172;
    output n5_adj_173;
    output n4_adj_174;
    output n7_adj_175;
    input n82;
    input n84;
    output n6_adj_176;
    output n9_adj_177;
    output n3_adj_178;
    output n8_adj_179;
    output n23_adj_180;
    output n7_adj_181;
    output n2_adj_182;
    output n5_adj_183;
    input n79;
    input n81_adj_184;
    output n9_adj_185;
    input n76;
    input n78_adj_186;
    output n4_adj_187;
    output n11_adj_188;
    output n10_adj_189;
    output n7_adj_190;
    output n6_adj_191;
    output n31_adj_192;
    output n9_adj_193;
    output n21_adj_194;
    output n20_adj_195;
    output n8_adj_196;
    output \d_out_11__N_1819[10] ;
    output n11_adj_197;
    output n13_adj_198;
    output n12_adj_199;
    output n30_adj_200;
    output n10_adj_201;
    output n13_adj_202;
    output \d_out_11__N_1819[11] ;
    output n8_adj_203;
    output n12_adj_204;
    output n15_adj_205;
    output n15_adj_206;
    output n14_adj_207;
    output n14_adj_208;
    output n17_adj_209;
    output n16_adj_210;
    output n19_adj_211;
    output n17_adj_212;
    output n18_adj_213;
    output n16_adj_214;
    output n21_adj_215;
    output n20_adj_216;
    output n19_adj_217;
    output n23_adj_218;
    output n22_adj_219;
    output n25_adj_220;
    output n18_adj_221;
    output n21_adj_222;
    output n20_adj_223;
    output \d_out_11__N_1819[8] ;
    output n24_adj_224;
    output n27_adj_225;
    output n23_adj_226;
    output \d_out_11__N_1819[9] ;
    output n22_adj_227;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(89[6:21])
    
    wire clk_80mhz_enable_141, clk_80mhz_enable_64, d_clk_tmp, n12602, 
        v_comb;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    
    wire n64_c, n132, clk_80mhz_enable_161, n65_c, n133, n18153, 
        n18157, n18156;
    wire [71:0]d10;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(47[26:29])
    
    wire n18166, n17821, n18165, n18169, n17810, n18168, n18172, 
        n18171, n18175, n18174, n17802, n18178, d_clk_tmp_N_1831, 
        n18177, n18181, n18180, n18187, n18186, n66, n134, clk_80mhz_enable_211, 
        clk_80mhz_enable_261, clk_80mhz_enable_311, clk_80mhz_enable_361, 
        clk_80mhz_enable_411, clk_80mhz_enable_461, clk_80mhz_enable_511, 
        clk_80mhz_enable_561, clk_80mhz_enable_611, clk_80mhz_enable_661, 
        clk_80mhz_enable_711;
    wire [71:0]d10_71__N_1747;
    
    wire n63, n12618, n67, n135, n136, n137, n131, n31_adj_2624, 
        n131_adj_2627, n132_adj_2633, n133_adj_2637, n134_adj_2640, 
        n135_adj_2642, n136_adj_2647, n17274, n17760, n17738, n17730, 
        n18269, n17756, n17734, n17617, n17633, n17637, n17635, 
        n18154;
    
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3JX d_clk_tmp_65 (.D(n12602), .CK(clk_80mhz), .PD(clk_80mhz_enable_141), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(clk_80mhz), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_64), 
            .CK(clk_80mhz), .Q(CIC1_outSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_141), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(n132), .Z(d_out_11__N_1819[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26_adj_115)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_64), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_116)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35_adj_117)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(n133), .Z(d_out_11__N_1819[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    LUT4 shift_right_31_i210_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[69] ), 
         .C(\d10[68] ), .Z(n18153)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[65] ), 
         .C(\d10[66] ), .Z(n18157)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[68] ), 
         .C(\d10[67] ), .Z(n18156)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 i6692_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n18166)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6692_then_3_lut.init = 16'he4e4;
    LUT4 i6692_else_3_lut (.A(n17821), .B(\CICGain[1] ), .C(d10[59]), 
         .Z(n18165)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6692_else_3_lut.init = 16'he2e2;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 i6650_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n18169)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6650_then_3_lut.init = 16'he4e4;
    LUT4 i6650_else_3_lut (.A(n17810), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n18168)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6650_else_3_lut.init = 16'he2e2;
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    LUT4 shift_right_31_i212_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(\d10[68] ), 
         .C(\d10[70] ), .Z(n18172)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_3_lut (.A(\d10[71] ), .B(\CICGain[1] ), 
         .C(\d10[69] ), .Z(n18171)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(\d10[67] ), .C(\d10[69] ), 
         .Z(n18175)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\d10[70] ), .B(\CICGain[1] ), .C(\d10[68] ), 
         .Z(n18174)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    LUT4 shift_right_31_i212_3_lut_4_lut_then_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[68]), .D(n17802), .Z(n18178)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((D)+!B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_then_4_lut.init = 16'hf791;
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_118)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34_adj_119)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    LUT4 shift_right_31_i212_3_lut_4_lut_else_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[68]), .D(n17802), .Z(n18177)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (D))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_else_4_lut.init = 16'he680;
    LUT4 i11_3_lut_4_lut_then_3_lut_adj_28 (.A(\CICGain[1] ), .B(d10[67]), 
         .C(d10[69]), .Z(n18181)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_then_3_lut_adj_28.init = 16'hd8d8;
    LUT4 shift_right_31_i62_rep_60_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n17821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i62_rep_60_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_29 (.A(d10[70]), .B(\CICGain[1] ), 
         .C(d10[68]), .Z(n18180)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_else_3_lut_adj_29.init = 16'he2e2;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37_adj_120)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_121)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_122)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36_adj_123)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 i6674_then_3_lut (.A(\CICGain[1] ), .B(d10[68]), .C(d10[66]), 
         .Z(n18187)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6674_then_3_lut.init = 16'he4e4;
    LUT4 i6674_else_3_lut (.A(n17802), .B(\CICGain[1] ), .C(d10[67]), 
         .Z(n18186)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6674_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(n134), .Z(d_out_11__N_1819[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_261), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_261), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_711), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1819[2]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1819[3]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1819[4]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1819[5]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1819[6]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1819[7]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1819[8]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1819[10]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1819[11]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    FD1S3IX count__i2 (.D(n87_adj_228[2]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_228[3]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_228[4]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_228[5]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_228[6]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_228[7]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_228[8]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_228[9]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_228[10]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(d_clk_tmp_N_1831), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_228[12]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_228[13]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_228[14]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_228[15]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n87_adj_228[1]), .CK(clk_80mhz), .CD(n12618), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(n135), .Z(d_out_11__N_1819[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[67]), .D(n136), .Z(d_out_11__N_1819[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i209_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[68]), .D(n137), .Z(d_out_11__N_1819[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i209_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_125), .D(n131), .Z(\d_out_11__N_1819[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11_adj_126)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10_adj_127)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17821), .D(d10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 i3134_2_lut (.A(n87_adj_228[0]), .B(n31_adj_2624), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(86[13] 89[16])
    defparam i3134_2_lut.init = 16'hbbbb;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_128)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_129)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_30 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(n131_adj_2627), .Z(d_out_11__N_1819[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_30.init = 16'hfe10;
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_130)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_131)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31_adj_132)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30_adj_133)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_31 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(n132_adj_2633), .Z(\d_out_11__N_1819[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_31.init = 16'hfe10;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_134)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_32 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(n133_adj_2637), .Z(\d_out_11__N_1819[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_32.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_33 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_135), .D(n134_adj_2640), .Z(\d_out_11__N_1819[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_33.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_34 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[66] ), .D(n135_adj_2642), .Z(\d_out_11__N_1819[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_34.init = 16'hfe10;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_136)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_137)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_35 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_135), .D(\d10[64] ), .Z(n136_adj_2647)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_35.init = 16'hf960;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15_adj_138)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_36 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(\d10[62] ), .Z(n134_adj_2640)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_36.init = 16'hf960;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_37 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(\d10[63] ), .Z(n135_adj_2642)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_37.init = 16'hf960;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_38 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17784), .D(\d10[60] ), .Z(n132_adj_2633)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_38.init = 16'hf960;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14_adj_139)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_140)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_39 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_125), .D(\d10[61] ), .Z(n133_adj_2637)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_39.init = 16'hf960;
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17805), .D(\d10[59] ), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 i6587_4_lut_rep_185 (.A(n17274), .B(n17760), .C(n17738), .D(n17730), 
         .Z(n18269)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(74[11:40])
    defparam i6587_4_lut_rep_185.init = 16'h4000;
    LUT4 shift_right_31_i137_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(d10[65]), .Z(n137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_141)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_40 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17810), .D(d10[59]), .Z(n131_adj_2627)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_40.init = 16'hf960;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5_adj_142)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4_adj_143)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i67_rep_66_3_lut (.A(d10[66]), .B(d10[67]), .C(\CICGain[0] ), 
         .Z(n67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i67_rep_66_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_41 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[67] ), .D(n136_adj_2647), .Z(\d_out_11__N_1819[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_41.init = 16'hfe10;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33_adj_144)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6_adj_145)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19_adj_146)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27_adj_147)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26_adj_148)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_196 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_511)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_196.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29_adj_149)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_191 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_261)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_191.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_190 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_211)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_190.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_195 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_461)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_195.GSR = "ENABLED";
    LUT4 i6587_4_lut_rep_186 (.A(n17274), .B(n17760), .C(n17738), .D(n17730), 
         .Z(clk_80mhz_enable_141)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(74[11:40])
    defparam i6587_4_lut_rep_186.init = 16'h4000;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22_adj_150)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_189 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_161)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_189.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_188 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_64)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_188.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28_adj_151)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 i6587_4_lut (.A(n17274), .B(n17760), .C(n17738), .D(n17730), 
         .Z(d_clk_tmp_N_1831)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(74[11:40])
    defparam i6587_4_lut.init = 16'h4000;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18_adj_152)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 i6547_4_lut (.A(n17756), .B(count[5]), .C(n17734), .D(count[9]), 
         .Z(n17760)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6547_4_lut.init = 16'h8000;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31_adj_153)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_154)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_155)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_156)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33_adj_157)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25_adj_158)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 mux_1252_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i2_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32_adj_159)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24_adj_160)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 i2865_2_lut (.A(n31_adj_2624), .B(d_clk_tmp), .Z(n12602)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam i2865_2_lut.init = 16'h8888;
    LUT4 mux_1252_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i3_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35_adj_161)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_162)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 i6526_2_lut (.A(count[2]), .B(count[4]), .Z(n17738)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6526_2_lut.init = 16'h8888;
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34_adj_163)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_164)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_165)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 mux_1252_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i4_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_166)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 mux_1252_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1252_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1252_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i7_3_lut.init = 16'hcaca;
    LUT4 i6518_2_lut (.A(count[8]), .B(count[3]), .Z(n17730)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6518_2_lut.init = 16'h8888;
    LUT4 i6543_3_lut (.A(count[6]), .B(count[7]), .C(count[10]), .Z(n17756)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i6543_3_lut.init = 16'h8080;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37_adj_167)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_168)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 mux_1252_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1252_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i9_3_lut.init = 16'hcaca;
    LUT4 i6522_2_lut (.A(count[0]), .B(count[1]), .Z(n17734)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6522_2_lut.init = 16'h8888;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36_adj_169)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 mux_1252_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i10_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(count[12]), .B(count[11]), .C(n17617), .D(count[15]), 
         .Z(n17274)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 mux_1252_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1252_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i12_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_170)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 mux_1252_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i13_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i70_rep_41_3_lut (.A(d10[69]), .B(d10[70]), .C(\CICGain[0] ), 
         .Z(n17802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i70_rep_41_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17617)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_171)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_172)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_173)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_200 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_711)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_200.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_42 (.A(n17633), .B(n17274), .C(n17637), .D(n17635), 
         .Z(n31_adj_2624)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_42.init = 16'hfffe;
    FD1S3AX v_comb_66_rep_199 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_661)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_199.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_198 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_611)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_198.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17633)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_43 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17637)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_43.init = 16'hfffe;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_174)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_44 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17635)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_44.init = 16'hfffe;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7_adj_175)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 mux_1252_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i14_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6_adj_176)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_177)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3_adj_178)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 i6592_2_lut (.A(n31_adj_2624), .B(n18269), .Z(n12618)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam i6592_2_lut.init = 16'hdddd;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_179)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_180)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_193 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_361)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_193.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7_adj_181)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2_adj_182)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 i3192_2_lut (.A(n87_adj_228[11]), .B(n31_adj_2624), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(86[13] 89[16])
    defparam i3192_2_lut.init = 16'hbbbb;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5_adj_183)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 mux_1252_i15_3_lut (.A(n79), .B(n81_adj_184), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i15_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_185)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    PFUMX i6718 (.BLUT(n18186), .ALUT(n18187), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[9]));
    LUT4 mux_1252_i16_3_lut (.A(n76), .B(n78_adj_186), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1252_i16_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4_adj_187)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_188)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    PFUMX i6714 (.BLUT(n18180), .ALUT(n18181), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[10]));
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_189)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_190)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_191)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    PFUMX i6712 (.BLUT(n18177), .ALUT(n18178), .C0(d10[71]), .Z(d_out_11__N_1819[11]));
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_192)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_193)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21_adj_194)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20_adj_195)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_196)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    PFUMX i6710 (.BLUT(n18174), .ALUT(n18175), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[10] ));
    LUT4 shift_right_31_i61_rep_49_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n17810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i61_rep_49_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11_adj_197)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13_adj_198)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12_adj_199)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30_adj_200)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_201)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_202)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    PFUMX i6708 (.BLUT(n18171), .ALUT(n18172), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[11] ));
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_203)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_204)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_205)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15_adj_206)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14_adj_207)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_208)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    PFUMX i6706 (.BLUT(n18168), .ALUT(n18169), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_209)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_210)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19_adj_211)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17_adj_212)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_213)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    PFUMX i6704 (.BLUT(n18165), .ALUT(n18166), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16_adj_214)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_215)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_216)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_217)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23_adj_218)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_192 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_311)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_192.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_219)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25_adj_220)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_221)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i210_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[66] ), 
         .C(\d10[67] ), .Z(n18154)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_222)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20_adj_223)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_197 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_561)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_197.GSR = "ENABLED";
    PFUMX i6698 (.BLUT(n18156), .ALUT(n18157), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[8] ));
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24_adj_224)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27_adj_225)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23_adj_226)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_194 (.D(clk_80mhz_enable_141), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_411)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=181, LSE_RLINE=187 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_194.GSR = "ENABLED";
    PFUMX i6696 (.BLUT(n18153), .ALUT(n18154), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[9] ));
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22_adj_227)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (clk_80mhz, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_80mhz;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_4_inv, rom_addr0_r_3_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, rom_dout_2_inv, rom_dout_1_inv, co0_1, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_4_inv, rom_dout_3_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_6_inv, rom_dout_5_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_8_inv, rom_dout_7_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_10_inv, rom_dout_9_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_12_inv, rom_dout_11_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_15_inv, 
        rom_dout_14_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_17_inv, 
        rom_dout_16_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_19_inv, 
        rom_dout_18_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_21_inv, 
        rom_dout_20_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_23_inv, 
        rom_dout_22_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_25_inv, 
        rom_dout_24_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    CCU2C neg_rom_addr0_r_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(702[11] 704[71])
    defparam neg_rom_addr0_r_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_0.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
          .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(710[11] 713[42])
    defparam neg_rom_addr0_r_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
          .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(719[11] 722[42])
    defparam neg_rom_addr0_r_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(728[11] 730[73])
    defparam neg_rom_addr0_r_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_3.INJECT1_1 = "NO";
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    CCU2C neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
          .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(874[11] 877[43])
    defparam neg_rom_dout_s_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
          .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(883[11] 886[43])
    defparam neg_rom_dout_s_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_6_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
          .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(892[11] 895[41])
    defparam neg_rom_dout_s_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_8_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
          .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(901[11] 904[41])
    defparam neg_rom_dout_s_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_10_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
          .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(910[11] 913[42])
    defparam neg_rom_dout_s_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_12_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5), .S0(rom_dout_s_n_11), .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(919[11] 922[42])
    defparam neg_rom_dout_s_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_6.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_13_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(936[11] 938[72])
    defparam neg_rom_dout_c_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_0.INJECT1_1 = "NO";
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    CCU2C neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_15_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
          .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(944[11] 947[43])
    defparam neg_rom_dout_c_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_17_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
          .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(953[11] 956[43])
    defparam neg_rom_dout_c_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_19_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
          .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(962[11] 965[43])
    defparam neg_rom_dout_c_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_21_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
          .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(971[11] 974[43])
    defparam neg_rom_dout_c_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_23_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
          .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(980[11] 983[44])
    defparam neg_rom_dout_c_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_25_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5_1), .S0(rom_dout_c_n_11), .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(989[11] 992[44])
    defparam neg_rom_dout_c_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_6.INJECT1_1 = "NO";
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(151[8] 158[2])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    CCU2C neg_rom_dout_s_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=158 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/SinCos/SinCos.v(866[11] 868[72])
    defparam neg_rom_dout_s_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_0.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PLL
//

module PLL (clk_25mhz_c, clk_80mhz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_25mhz_c;
    output clk_80mhz;
    input GND_net;
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(68[8:17])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    
    EHXPLLL PLLInst_0 (.CLKI(clk_25mhz_c), .CLKFB(clk_80mhz), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .PHASELOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .CLKOP(clk_80mhz)) /* synthesis FREQUENCY_PIN_CLKOP="83.333333", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="5", LPF_RESISTOR="16", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=145, LSE_RLINE=148 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(145[5] 148[2])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.CLKOP_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.PLL_LOCK_DELAY = 200;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.REFIN_RESET = "DISABLED";
    defparam PLLInst_0.SYNC_ENABLE = "DISABLED";
    defparam PLLInst_0.INT_LOCK_STICKY = "ENABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module nco_sig
//

module nco_sig (\phase_accum[63] , sinGen_c) /* synthesis syn_module_defined=1 */ ;
    input \phase_accum[63] ;
    output sinGen_c;
    
    
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/NCO.v(32[18:56])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096)_U1 
//

module \CIC(width=72,decimation_ratio=4096)_U1  (d_d8, n3, d_tmp, clk_80mhz, 
            d5, d_d_tmp, d2, d2_71__N_490, d3, d3_71__N_562, d4, 
            d4_71__N_634, d5_71__N_706, d6, d6_71__N_1459, d_d6, d7, 
            d7_71__N_1531, d_d7, d8, d8_71__N_1603, d9, d9_71__N_1675, 
            d_d9, CIC1_outCos, d1, d1_71__N_418, n15, count, n28, 
            n14, n2, n87_adj_114, n17, n3_adj_1, n9, n2_adj_2, 
            n5, n8, n4, n7, n23, n22, n2_adj_3, n25, n5_adj_4, 
            n4_adj_5, \CICGain[1] , \d10[60] , n17784, \d10[59] , 
            n24, n27, n26, n29, n28_adj_6, n31, n30, n7_adj_7, 
            n33, n6, n6_adj_8, n11, n10, n32, n9_adj_9, n8_adj_10, 
            n35, n34, n17805, \d10[62] , \d10[63] , \CICGain[0] , 
            n63_adj_11, n37, n29_adj_12, n5_adj_13, n36_adj_14, n16, 
            n13, n12, n15_adj_15, n14_adj_16, n17_adj_17, n16_adj_18, 
            n19, n18, n21, n20, \d10[61] , \d10[64] , \d10[65] , 
            \d10[66] , \d10[67] , \d10[68] , \d10[69] , \d10[70] , 
            \d10[71] , \d_out_11__N_1819[2] , \d_out_11__N_1819[3] , \d_out_11__N_1819[4] , 
            \d_out_11__N_1819[5] , \d_out_11__N_1819[6] , \d_out_11__N_1819[7] , 
            \d_out_11__N_1819[8] , \d_out_11__N_1819[9] , \d_out_11__N_1819[10] , 
            \d_out_11__N_1819[11] , n19_adj_19, n11_adj_20, n33_adj_21, 
            n32_adj_22, n35_adj_23, n10_adj_24, n13_adj_25, n12_adj_26, 
            n15_adj_27, n14_adj_28, n17_adj_29, n16_adj_30, n19_adj_31, 
            n18_adj_32, n21_adj_33, n20_adj_34, n23_adj_35, n22_adj_36, 
            n25_adj_37, n24_adj_38, n3_adj_39, n27_adj_40, n26_adj_41, 
            n2_adj_42, n5_adj_43, n29_adj_44, n28_adj_45, n4_adj_46, 
            n7_adj_47, n31_adj_48, n30_adj_49, n6_adj_50, n9_adj_51, 
            n33_adj_52, n32_adj_53, n8_adj_54, n11_adj_55, n35_adj_56, 
            n34_adj_57, n4_adj_58, n10_adj_59, n13_adj_60, n34_adj_61, 
            n23_adj_62, n22_adj_63, n27_adj_64, n26_adj_65, n37_adj_66, 
            n36_adj_67, n12_adj_68, n18_adj_69, n21_adj_70, n64, n7_adj_71, 
            n65, n20_adj_72, n18_adj_73, n23_adj_74, n22_adj_75, n21_adj_76, 
            n6_adj_77, n25_adj_78, n24_adj_79, n66_adj_80, n9_adj_81, 
            n8_adj_82, n27_adj_83, n11_adj_84, n10_adj_85, n26_adj_86, 
            n29_adj_87, n28_adj_88, n31_adj_89, n30_adj_90, n13_adj_91, 
            n33_adj_92, n32_adj_93, n12_adj_94, n35_adj_95, n15_adj_96, 
            n34_adj_97, n31_adj_98, n30_adj_99, n37_adj_100, n14_adj_101, 
            n36_adj_102, n20_adj_103, n17_adj_104, n16_adj_105, n19_adj_106, 
            n118, n120, cout, n115, n117, n112, n114, n109, 
            n111, n106, n108, n37_adj_107, n36_adj_108, n103, n105, 
            n100, n102, n97, n99, n94, n96, n91, n93, n25_adj_109, 
            n88, n90, n24_adj_110, n85, n87, n82, n84, n79, 
            n81_adj_111, n76, n78_adj_112, n3_adj_113) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_d8;
    output n3;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d_d7;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output [11:0]CIC1_outCos;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output n15;
    output [15:0]count;
    output n28;
    output n14;
    output n2;
    input [15:0]n87_adj_114;
    output n17;
    output n3_adj_1;
    output n9;
    output n2_adj_2;
    output n5;
    output n8;
    output n4;
    output n7;
    output n23;
    output n22;
    output n2_adj_3;
    output n25;
    output n5_adj_4;
    output n4_adj_5;
    input \CICGain[1] ;
    output \d10[60] ;
    output n17784;
    output \d10[59] ;
    output n24;
    output n27;
    output n26;
    output n29;
    output n28_adj_6;
    output n31;
    output n30;
    output n7_adj_7;
    output n33;
    output n6;
    output n6_adj_8;
    output n11;
    output n10;
    output n32;
    output n9_adj_9;
    output n8_adj_10;
    output n35;
    output n34;
    output n17805;
    output \d10[62] ;
    output \d10[63] ;
    input \CICGain[0] ;
    output n63_adj_11;
    output n37;
    output n29_adj_12;
    output n5_adj_13;
    output n36_adj_14;
    output n16;
    output n13;
    output n12;
    output n15_adj_15;
    output n14_adj_16;
    output n17_adj_17;
    output n16_adj_18;
    output n19;
    output n18;
    output n21;
    output n20;
    output \d10[61] ;
    output \d10[64] ;
    output \d10[65] ;
    output \d10[66] ;
    output \d10[67] ;
    output \d10[68] ;
    output \d10[69] ;
    output \d10[70] ;
    output \d10[71] ;
    input \d_out_11__N_1819[2] ;
    input \d_out_11__N_1819[3] ;
    input \d_out_11__N_1819[4] ;
    input \d_out_11__N_1819[5] ;
    input \d_out_11__N_1819[6] ;
    input \d_out_11__N_1819[7] ;
    input \d_out_11__N_1819[8] ;
    input \d_out_11__N_1819[9] ;
    input \d_out_11__N_1819[10] ;
    input \d_out_11__N_1819[11] ;
    output n19_adj_19;
    output n11_adj_20;
    output n33_adj_21;
    output n32_adj_22;
    output n35_adj_23;
    output n10_adj_24;
    output n13_adj_25;
    output n12_adj_26;
    output n15_adj_27;
    output n14_adj_28;
    output n17_adj_29;
    output n16_adj_30;
    output n19_adj_31;
    output n18_adj_32;
    output n21_adj_33;
    output n20_adj_34;
    output n23_adj_35;
    output n22_adj_36;
    output n25_adj_37;
    output n24_adj_38;
    output n3_adj_39;
    output n27_adj_40;
    output n26_adj_41;
    output n2_adj_42;
    output n5_adj_43;
    output n29_adj_44;
    output n28_adj_45;
    output n4_adj_46;
    output n7_adj_47;
    output n31_adj_48;
    output n30_adj_49;
    output n6_adj_50;
    output n9_adj_51;
    output n33_adj_52;
    output n32_adj_53;
    output n8_adj_54;
    output n11_adj_55;
    output n35_adj_56;
    output n34_adj_57;
    output n4_adj_58;
    output n10_adj_59;
    output n13_adj_60;
    output n34_adj_61;
    output n23_adj_62;
    output n22_adj_63;
    output n27_adj_64;
    output n26_adj_65;
    output n37_adj_66;
    output n36_adj_67;
    output n12_adj_68;
    output n18_adj_69;
    output n21_adj_70;
    output n64;
    output n7_adj_71;
    output n65;
    output n20_adj_72;
    output n18_adj_73;
    output n23_adj_74;
    output n22_adj_75;
    output n21_adj_76;
    output n6_adj_77;
    output n25_adj_78;
    output n24_adj_79;
    output n66_adj_80;
    output n9_adj_81;
    output n8_adj_82;
    output n27_adj_83;
    output n11_adj_84;
    output n10_adj_85;
    output n26_adj_86;
    output n29_adj_87;
    output n28_adj_88;
    output n31_adj_89;
    output n30_adj_90;
    output n13_adj_91;
    output n33_adj_92;
    output n32_adj_93;
    output n12_adj_94;
    output n35_adj_95;
    output n15_adj_96;
    output n34_adj_97;
    output n31_adj_98;
    output n30_adj_99;
    output n37_adj_100;
    output n14_adj_101;
    output n36_adj_102;
    output n20_adj_103;
    output n17_adj_104;
    output n16_adj_105;
    output n19_adj_106;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    input n109;
    input n111;
    input n106;
    input n108;
    output n37_adj_107;
    output n36_adj_108;
    input n103;
    input n105;
    input n100;
    input n102;
    input n97;
    input n99;
    input n94;
    input n96;
    input n91;
    input n93;
    output n25_adj_109;
    input n88;
    input n90;
    output n24_adj_110;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81_adj_111;
    input n76;
    input n78_adj_112;
    output n3_adj_113;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(72[6:15])
    
    wire clk_80mhz_enable_758, clk_80mhz_enable_798, v_comb;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    
    wire n31_c, n18285, n12630;
    wire [71:0]d10;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(47[26:29])
    
    wire n18160, n18159, n18184, n18183, n17266, n17758, n17728, 
        n17720, count_15__N_1458, n17748, clk_80mhz_enable_910, clk_80mhz_enable_960, 
        clk_80mhz_enable_1010, clk_80mhz_enable_1060, clk_80mhz_enable_1110, 
        clk_80mhz_enable_1160, clk_80mhz_enable_1210, clk_80mhz_enable_1260, 
        clk_80mhz_enable_1310, clk_80mhz_enable_1360, clk_80mhz_enable_1410, 
        clk_80mhz_enable_1460;
    wire [71:0]d10_71__N_1747;
    
    wire n17663, n17653, n17657, n17655;
    
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_798), 
            .CK(clk_80mhz), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_758), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 i6619_2_lut (.A(n31_c), .B(n18285), .Z(n12630)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam i6619_2_lut.init = 16'hdddd;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 i3193_2_lut (.A(n87_adj_114[11]), .B(n31_c), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(86[13] 89[16])
    defparam i3193_2_lut.init = 16'hbbbb;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_1)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2_adj_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5_adj_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4_adj_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 i6666_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n18160)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6666_then_3_lut.init = 16'he4e4;
    LUT4 i6666_else_3_lut (.A(n17784), .B(\CICGain[1] ), .C(\d10[59] ), 
         .Z(n18159)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6666_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28_adj_6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7_adj_7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6_adj_8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 i6680_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n18184)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6680_then_3_lut.init = 16'he4e4;
    LUT4 i6680_else_3_lut (.A(n17805), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n18183)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6680_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63_adj_11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5_adj_13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36_adj_14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15_adj_15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14_adj_16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17_adj_17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16_adj_18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 i6581_4_lut (.A(n17266), .B(n17758), .C(n17728), .D(n17720), 
         .Z(count_15__N_1458)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(74[11:40])
    defparam i6581_4_lut.init = 16'h4000;
    LUT4 i6545_4_lut (.A(count[0]), .B(n17748), .C(count[6]), .D(count[10]), 
         .Z(n17758)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6545_4_lut.init = 16'h8000;
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_910), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_910), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_960), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_1010), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_1010), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_1010), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_1060), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_1060), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_1110), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_1110), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_1110), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_1110), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_1110), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_1110), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_1110), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_1160), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_1210), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_1210), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_1260), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_1260), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_1310), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_1360), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_1360), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_1410), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_1410), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_1460), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1819[2] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1819[3] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1819[4] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1819[5] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1819[6] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1819[7] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1819[8] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(\d_out_11__N_1819[9] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1819[10] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1819[11] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 i6516_2_lut (.A(count[2]), .B(count[4]), .Z(n17728)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6516_2_lut.init = 16'h8888;
    LUT4 i6508_2_lut (.A(count[7]), .B(count[3]), .Z(n17720)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6508_2_lut.init = 16'h8888;
    LUT4 i6535_4_lut (.A(count[5]), .B(count[1]), .C(count[9]), .D(count[8]), 
         .Z(n17748)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6535_4_lut.init = 16'h8000;
    FD1S3IX count__i2 (.D(n87_adj_114[2]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_114[3]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_114[4]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_114[5]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_114[6]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_114[7]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_114[8]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_114[9]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_114[10]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(count_15__N_1458), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_114[12]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_114[13]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_114[14]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_114[15]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(count[12]), .B(count[11]), .C(n17663), .D(count[15]), 
         .Z(n17266)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17663)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35_adj_23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10_adj_24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15_adj_27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14_adj_28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19_adj_31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18_adj_32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21_adj_33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20_adj_34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22_adj_36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25_adj_37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24_adj_38)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_39)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27_adj_40)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26_adj_41)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_42)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_43)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29_adj_44)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28_adj_45)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_46)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7_adj_47)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31_adj_48)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_49)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6_adj_50)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_51)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33_adj_52)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32_adj_53)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_54)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_55)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35_adj_56)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34_adj_57)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4_adj_58)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_59)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13_adj_60)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 i6581_4_lut_rep_201 (.A(n17266), .B(n17758), .C(n17728), .D(n17720), 
         .Z(n18285)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(74[11:40])
    defparam i6581_4_lut_rep_201.init = 16'h4000;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34_adj_61)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 i6581_4_lut_rep_202 (.A(n17266), .B(n17758), .C(n17728), .D(n17720), 
         .Z(clk_80mhz_enable_758)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(74[11:40])
    defparam i6581_4_lut_rep_202.init = 16'h4000;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23_adj_62)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22_adj_63)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_64)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_65)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37_adj_66)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_67)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12_adj_68)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_44_3_lut (.A(\d10[60] ), .B(\d10[61] ), 
         .C(\CICGain[0] ), .Z(n17805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i61_rep_44_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_69)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_211 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1210)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_211.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_210 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1160)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_210.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_70)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_209 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1110)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_209.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_208 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1060)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_208.GSR = "ENABLED";
    LUT4 shift_right_31_i64_3_lut (.A(\d10[63] ), .B(\d10[64] ), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_71)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i65_3_lut (.A(\d10[64] ), .B(\d10[65] ), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20_adj_72)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 i3136_2_lut (.A(n87_adj_114[0]), .B(n31_c), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(86[13] 89[16])
    defparam i3136_2_lut.init = 16'hbbbb;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_73)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_25 (.A(n17653), .B(n17266), .C(n17657), .D(n17655), 
         .Z(n31_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_25.init = 16'hfffe;
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17653)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_26 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17657)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_26.init = 16'hfffe;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23_adj_74)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22_adj_75)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_27 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17655)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_27.init = 16'hfffe;
    FD1S3AX v_comb_66_rep_207 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1010)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_207.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_206 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_960)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_206.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_76)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_77)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25_adj_78)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24_adj_79)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66_adj_80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_81)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_82)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27_adj_83)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11_adj_84)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_85)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_86)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_87)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_88)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31_adj_89)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30_adj_90)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_91)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33_adj_92)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32_adj_93)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_94)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_95)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_96)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_97)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_98)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_205 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_910)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_205.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_204 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_798)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_204.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30_adj_99)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37_adj_100)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_101)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36_adj_102)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_103)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_104)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_105)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19_adj_106)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 mux_1250_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i5_3_lut.init = 16'hcaca;
    PFUMX i6716 (.BLUT(n18183), .ALUT(n18184), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    LUT4 mux_1250_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i6_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_107)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_108)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 mux_1250_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i8_3_lut.init = 16'hcaca;
    FD1S3IX count__i1 (.D(n87_adj_114[1]), .CK(clk_80mhz), .CD(n12630), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 mux_1250_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i11_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_109)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 mux_1250_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i12_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_110)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 mux_1250_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i15_3_lut (.A(n79), .B(n81_adj_111), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i16_3_lut (.A(n76), .B(n78_adj_112), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(115[18:27])
    defparam mux_1250_i16_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3_adj_113)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_216 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1460)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_216.GSR = "ENABLED";
    PFUMX i6700 (.BLUT(n18159), .ALUT(n18160), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    FD1S3AX v_comb_66_rep_215 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1410)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_215.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_214 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1360)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_214.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_213 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1310)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_213.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_212 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1260)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_212.GSR = "ENABLED";
    LUT4 shift_right_31_i62_rep_23_3_lut (.A(\d10[61] ), .B(\d10[62] ), 
         .C(\CICGain[0] ), .Z(n17784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/CIC.v(119[20:47])
    defparam shift_right_31_i62_rep_23_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (\d_out_d_11__N_1892[17] , CIC1_out_clkSin, CIC1_outSin, 
            CIC1_outCos, \DataInReg_11__N_1856[0] , \d_out_d_11__N_1890[17] , 
            \d_out_d_11__N_1888[17] , \d_out_d_11__N_1886[17] , \d_out_d_11__N_1884[17] , 
            \d_out_d_11__N_1882[17] , \d_out_d_11__N_1880[17] , d_out_d_11__N_1879, 
            \d_out_d_11__N_1878[17] , d_out_d_11__N_1877, \d_out_d_11__N_1876[17] , 
            d_out_d_11__N_1875, \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , 
            \DataInReg_11__N_1856[3] , \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , 
            \DataInReg_11__N_1856[6] , \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] , 
            \DemodOut[9] , \ISquare[31] , n209, \d_out_d_11__N_2335[17] , 
            \d_out_d_11__N_2353[17] , \d_out_d_11__N_1874[17] , d_out_d_11__N_1873, 
            VCC_net, GND_net, MultResult2, MultResult1) /* synthesis syn_module_defined=1 */ ;
    input \d_out_d_11__N_1892[17] ;
    input CIC1_out_clkSin;
    input [11:0]CIC1_outSin;
    input [11:0]CIC1_outCos;
    output \DataInReg_11__N_1856[0] ;
    input \d_out_d_11__N_1890[17] ;
    input \d_out_d_11__N_1888[17] ;
    input \d_out_d_11__N_1886[17] ;
    input \d_out_d_11__N_1884[17] ;
    input \d_out_d_11__N_1882[17] ;
    input \d_out_d_11__N_1880[17] ;
    output d_out_d_11__N_1879;
    input \d_out_d_11__N_1878[17] ;
    output d_out_d_11__N_1877;
    input \d_out_d_11__N_1876[17] ;
    output d_out_d_11__N_1875;
    output \DataInReg_11__N_1856[1] ;
    output \DataInReg_11__N_1856[2] ;
    output \DataInReg_11__N_1856[3] ;
    output \DataInReg_11__N_1856[4] ;
    output \DataInReg_11__N_1856[5] ;
    output \DataInReg_11__N_1856[6] ;
    output \DataInReg_11__N_1856[7] ;
    output \DataInReg_11__N_1856[8] ;
    output \DemodOut[9] ;
    input \ISquare[31] ;
    output n209;
    input \d_out_d_11__N_2335[17] ;
    input \d_out_d_11__N_2353[17] ;
    input \d_out_d_11__N_1874[17] ;
    output d_out_d_11__N_1873;
    input VCC_net;
    input GND_net;
    output [23:0]MultResult2;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(89[6:21])
    
    wire d_out_d_11__N_1891;
    wire [11:0]MultDataB;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(29[21:30])
    wire [11:0]MultDataC;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(33[21:30])
    wire [15:0]d_out_d;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(20[21:28])
    wire [17:0]d_out_d_11__N_1894;
    
    wire d_out_d_11__N_1889, d_out_d_11__N_1887, d_out_d_11__N_1885, d_out_d_11__N_1883, 
        d_out_d_11__N_1881;
    
    LUT4 d_out_d_11__I_10_1_lut (.A(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1891)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    FD1S3AX MultDataB_i0 (.D(CIC1_outSin[0]), .CK(CIC1_out_clkSin), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i0.GSR = "ENABLED";
    FD1S3AX MultDataC_i0 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), .Q(MultDataC[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i0.GSR = "ENABLED";
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i1.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    LUT4 d_out_d_11__I_9_1_lut (.A(\d_out_d_11__N_1890[17] ), .Z(d_out_d_11__N_1889)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(\d_out_d_11__N_1888[17] ), .Z(d_out_d_11__N_1887)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(\d_out_d_11__N_1886[17] ), .Z(d_out_d_11__N_1885)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(\d_out_d_11__N_1884[17] ), .Z(d_out_d_11__N_1883)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(\d_out_d_11__N_1882[17] ), .Z(d_out_d_11__N_1881)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_4_1_lut (.A(\d_out_d_11__N_1880[17] ), .Z(d_out_d_11__N_1879)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(\d_out_d_11__N_1878[17] ), .Z(d_out_d_11__N_1877)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_2_1_lut (.A(\d_out_d_11__N_1876[17] ), .Z(d_out_d_11__N_1875)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    FD1S3AX MultDataB_i1 (.D(CIC1_outSin[1]), .CK(CIC1_out_clkSin), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i1.GSR = "ENABLED";
    FD1S3AX MultDataB_i2 (.D(CIC1_outSin[2]), .CK(CIC1_out_clkSin), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i2.GSR = "ENABLED";
    FD1S3AX MultDataB_i3 (.D(CIC1_outSin[3]), .CK(CIC1_out_clkSin), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i3.GSR = "ENABLED";
    FD1S3AX MultDataB_i4 (.D(CIC1_outSin[4]), .CK(CIC1_out_clkSin), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i4.GSR = "ENABLED";
    FD1S3AX MultDataB_i5 (.D(CIC1_outSin[5]), .CK(CIC1_out_clkSin), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i5.GSR = "ENABLED";
    FD1S3AX MultDataB_i6 (.D(CIC1_outSin[6]), .CK(CIC1_out_clkSin), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i6.GSR = "ENABLED";
    FD1S3AX MultDataB_i7 (.D(CIC1_outSin[7]), .CK(CIC1_out_clkSin), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i7.GSR = "ENABLED";
    FD1S3AX MultDataB_i8 (.D(CIC1_outSin[8]), .CK(CIC1_out_clkSin), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i8.GSR = "ENABLED";
    FD1S3AX MultDataB_i9 (.D(CIC1_outSin[9]), .CK(CIC1_out_clkSin), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i9.GSR = "ENABLED";
    FD1S3AX MultDataB_i10 (.D(CIC1_outSin[10]), .CK(CIC1_out_clkSin), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i10.GSR = "ENABLED";
    FD1S3AX MultDataB_i11 (.D(CIC1_outSin[11]), .CK(CIC1_out_clkSin), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i11.GSR = "ENABLED";
    FD1S3AX MultDataC_i1 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), .Q(MultDataC[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i1.GSR = "ENABLED";
    FD1S3AX MultDataC_i2 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), .Q(MultDataC[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i2.GSR = "ENABLED";
    FD1S3AX MultDataC_i3 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), .Q(MultDataC[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i3.GSR = "ENABLED";
    FD1S3AX MultDataC_i4 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), .Q(MultDataC[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i4.GSR = "ENABLED";
    FD1S3AX MultDataC_i5 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), .Q(MultDataC[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i5.GSR = "ENABLED";
    FD1S3AX MultDataC_i6 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), .Q(MultDataC[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i6.GSR = "ENABLED";
    FD1S3AX MultDataC_i7 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), .Q(MultDataC[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i7.GSR = "ENABLED";
    FD1S3AX MultDataC_i8 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), .Q(MultDataC[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i8.GSR = "ENABLED";
    FD1S3AX MultDataC_i9 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), .Q(MultDataC[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i9.GSR = "ENABLED";
    FD1S3AX MultDataC_i10 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), .Q(MultDataC[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i10.GSR = "ENABLED";
    FD1S3AX MultDataC_i11 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), .Q(MultDataC[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i11.GSR = "ENABLED";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=222, LSE_RLINE=227 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i10.GSR = "ENABLED";
    LUT4 i1339_1_lut (.A(\ISquare[31] ), .Z(n209)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1339_1_lut.init = 16'h5555;
    LUT4 mux_82_i1_3_lut (.A(\d_out_d_11__N_2335[17] ), .B(\d_out_d_11__N_2353[17] ), 
         .C(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1894[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(60[11:28])
    defparam mux_82_i1_3_lut.init = 16'h3535;
    LUT4 d_out_d_11__I_1_1_lut (.A(\d_out_d_11__N_1874[17] ), .Z(d_out_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1891), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1889), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1887), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1885), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1883), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1881), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1879), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1877), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1875), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    Multiplier Multiplier2 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataC({MultDataC}), .MultResult2({MultResult2})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    Multiplier_U0 Multiplier1 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataB({MultDataB}), .MultResult1({MultResult1})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    
endmodule
//
// Verilog Description of module Multiplier
//

module Multiplier (CIC1_out_clkSin, VCC_net, GND_net, MultDataC, MultResult2) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataC;
    output [23:0]MultResult2;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(89[6:21])
    
    wire regb_b_1, Multiplier_0_mult_0_5_n1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, regb_b_3, Multiplier_0_mult_2_5_n1, Multiplier_0_pp_2_4, 
        regb_b_4, regb_b_5, Multiplier_0_mult_4_5_n1, Multiplier_0_pp_3_6, 
        regb_b_6, regb_b_7, Multiplier_0_mult_6_5_n1, Multiplier_0_pp_4_8, 
        regb_b_8, regb_b_9, Multiplier_0_mult_8_5_n1, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_10, 
        s_Multiplier_0_3_9, co_Multiplier_0_3_5, s_Multiplier_0_3_12, 
        s_Multiplier_0_3_11, co_Multiplier_0_3_6, s_Multiplier_0_3_14, 
        s_Multiplier_0_3_13, co_Multiplier_0_3_7, s_Multiplier_0_3_16, 
        s_Multiplier_0_3_15, co_Multiplier_0_3_8, s_Multiplier_0_3_18, 
        s_Multiplier_0_3_17, co_Multiplier_0_3_9, s_Multiplier_0_3_20, 
        s_Multiplier_0_3_19, co_Multiplier_0_3_10, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_21, s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, 
        co_t_Multiplier_0_4_2, co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, 
        co_t_Multiplier_0_4_5, co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, 
        co_t_Multiplier_0_4_8, mco, mco_1, mco_2, mco_3, mco_4, 
        Multiplier_0_mult_0_5_n2, mco_5, mco_6, mco_7, mco_8, mco_9, 
        Multiplier_0_mult_2_5_n2, mco_10, mco_11, mco_12, mco_13, 
        mco_14, Multiplier_0_mult_4_5_n2, mco_15, mco_16, mco_17, 
        mco_18, mco_19, Multiplier_0_mult_6_5_n2, mco_20, mco_21, 
        mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, Multiplier_0_mult_10_0_n1, 
        mco_25, mco_26, mco_27, mco_28, mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    FD1P3DX FF_98 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataC[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    CCU2C Multiplier_0_cin_lr_add_0 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(788[11] 790[76])
    defparam Multiplier_0_cin_lr_add_0.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_0.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_0.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_0_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(796[11] 798[79])
    defparam Multiplier_0_Cadd_0_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_0_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_0_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_0_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_2 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(804[11] 806[76])
    defparam Multiplier_0_cin_lr_add_2.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_2.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_2.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_2_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(812[11] 815[17])
    defparam Multiplier_0_Cadd_2_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_2_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_2_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_2_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_4 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(821[11] 823[76])
    defparam Multiplier_0_cin_lr_add_4.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_4.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_4.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_4_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(829[11] 832[17])
    defparam Multiplier_0_Cadd_4_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_4_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_4_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_4_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_6 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(838[11] 840[76])
    defparam Multiplier_0_cin_lr_add_6.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_6.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_6.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_6_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(846[11] 849[17])
    defparam Multiplier_0_Cadd_6_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_6_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_6_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_6_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_8 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(855[11] 857[76])
    defparam Multiplier_0_cin_lr_add_8.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_8.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_8.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_8.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_8_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(863[11] 866[17])
    defparam Multiplier_0_Cadd_8_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_8_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_8_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_8_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_10 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(872[11] 874[77])
    defparam Multiplier_0_cin_lr_add_10.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_10.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_10.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_10.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_10_6 (.A0(VCC_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(880[11] 883[17])
    defparam Multiplier_0_Cadd_10_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_10_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_10_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_10_6.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_0_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(Multiplier_0_pp_0_2), .B1(Multiplier_0_pp_1_2), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_0_1), .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(889[11] 892[36])
    defparam Cadd_Multiplier_0_0_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_0_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .B0(Multiplier_0_pp_1_3), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_4), .B1(Multiplier_0_pp_1_4), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_1), .COUT(co_Multiplier_0_0_2), 
          .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(898[11] 901[86])
    defparam Multiplier_0_add_0_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .B0(Multiplier_0_pp_1_5), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_6), .B1(Multiplier_0_pp_1_6), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_2), .COUT(co_Multiplier_0_0_3), 
          .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(907[11] 910[86])
    defparam Multiplier_0_add_0_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .B0(Multiplier_0_pp_1_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_8), .B1(Multiplier_0_pp_1_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_3), .COUT(co_Multiplier_0_0_4), 
          .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(916[11] 919[86])
    defparam Multiplier_0_add_0_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .B0(Multiplier_0_pp_1_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_10), .B1(Multiplier_0_pp_1_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_4), .COUT(co_Multiplier_0_0_5), 
          .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(925[11] 928[87])
    defparam Multiplier_0_add_0_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .B0(Multiplier_0_pp_1_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_12), .B1(Multiplier_0_pp_1_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_5), .COUT(co_Multiplier_0_0_6), 
          .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(934[11] 937[88])
    defparam Multiplier_0_add_0_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .B0(Multiplier_0_pp_1_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(Multiplier_0_pp_1_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_6), .COUT(co_Multiplier_0_0_7), 
          .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(943[11] 946[88])
    defparam Multiplier_0_add_0_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_8 (.A0(GND_net), .B0(Multiplier_0_pp_1_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
          .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(952[11] 955[62])
    defparam Multiplier_0_add_0_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_8.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_0_9 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(961[11] 964[24])
    defparam Cadd_Multiplier_0_0_9.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_9.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_9.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_0_9.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_1_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(Multiplier_0_pp_2_6), .B1(Multiplier_0_pp_3_6), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_1_1), .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(970[11] 973[36])
    defparam Cadd_Multiplier_0_1_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_1_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .B0(Multiplier_0_pp_3_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_8), .B1(Multiplier_0_pp_3_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_1), .COUT(co_Multiplier_0_1_2), 
          .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(979[11] 982[86])
    defparam Multiplier_0_add_1_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .B0(Multiplier_0_pp_3_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_10), .B1(Multiplier_0_pp_3_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_2), .COUT(co_Multiplier_0_1_3), 
          .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(988[11] 991[87])
    defparam Multiplier_0_add_1_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .B0(Multiplier_0_pp_3_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_12), .B1(Multiplier_0_pp_3_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_3), .COUT(co_Multiplier_0_1_4), 
          .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(997[11] 1000[88])
    defparam Multiplier_0_add_1_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .B0(Multiplier_0_pp_3_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_14), .B1(Multiplier_0_pp_3_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_4), .COUT(co_Multiplier_0_1_5), 
          .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1006[11] 1009[88])
    defparam Multiplier_0_add_1_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .B0(Multiplier_0_pp_3_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_16), .B1(Multiplier_0_pp_3_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_5), .COUT(co_Multiplier_0_1_6), 
          .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1015[11] 1018[88])
    defparam Multiplier_0_add_1_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .B0(Multiplier_0_pp_3_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(Multiplier_0_pp_3_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_6), .COUT(co_Multiplier_0_1_7), 
          .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1024[11] 1027[88])
    defparam Multiplier_0_add_1_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_8 (.A0(GND_net), .B0(Multiplier_0_pp_3_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
          .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1033[11] 1036[62])
    defparam Multiplier_0_add_1_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_8.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_1_9 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1042[11] 1045[24])
    defparam Cadd_Multiplier_0_1_9.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_9.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_9.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_1_9.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_2_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(Multiplier_0_pp_4_10), .B1(Multiplier_0_pp_5_10), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_2_1), .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1051[11] 1054[36])
    defparam Cadd_Multiplier_0_2_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_2_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_2_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_2_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .B0(Multiplier_0_pp_5_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_12), .B1(Multiplier_0_pp_5_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_1), .COUT(co_Multiplier_0_2_2), 
          .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1060[11] 1063[88])
    defparam Multiplier_0_add_2_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .B0(Multiplier_0_pp_5_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_14), .B1(Multiplier_0_pp_5_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_2), .COUT(co_Multiplier_0_2_3), 
          .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1069[11] 1072[88])
    defparam Multiplier_0_add_2_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .B0(Multiplier_0_pp_5_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_16), .B1(Multiplier_0_pp_5_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_3), .COUT(co_Multiplier_0_2_4), 
          .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1078[11] 1081[88])
    defparam Multiplier_0_add_2_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .B0(Multiplier_0_pp_5_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_18), .B1(Multiplier_0_pp_5_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_4), .COUT(co_Multiplier_0_2_5), 
          .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1087[11] 1090[88])
    defparam Multiplier_0_add_2_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .B0(Multiplier_0_pp_5_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_20), .B1(Multiplier_0_pp_5_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_5), .COUT(co_Multiplier_0_2_6), 
          .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1096[11] 1099[88])
    defparam Multiplier_0_add_2_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .B0(Multiplier_0_pp_5_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(Multiplier_0_pp_5_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_6), .COUT(co_Multiplier_0_2_7), 
          .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1105[11] 1108[88])
    defparam Multiplier_0_add_2_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_8 (.A0(GND_net), .B0(Multiplier_0_pp_5_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1114[11] 1117[43])
    defparam Multiplier_0_add_2_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_8.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_3_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(f_s_Multiplier_0_0_4), .B1(f_Multiplier_0_pp_2_4), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_3_1), .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1123[11] 1126[36])
    defparam Cadd_Multiplier_0_3_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_3_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .B0(f_Multiplier_0_pp_2_5), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_6), .B1(f_s_Multiplier_0_1_6), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_1), .COUT(co_Multiplier_0_3_2), 
          .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1132[11] 1135[86])
    defparam Multiplier_0_add_3_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .B0(f_s_Multiplier_0_1_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_8), .B1(f_s_Multiplier_0_1_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_2), .COUT(co_Multiplier_0_3_3), 
          .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1141[11] 1144[86])
    defparam Multiplier_0_add_3_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .B0(f_s_Multiplier_0_1_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_10), .B1(f_s_Multiplier_0_1_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_3), .COUT(co_Multiplier_0_3_4), 
          .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1150[11] 1153[87])
    defparam Multiplier_0_add_3_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .B0(f_s_Multiplier_0_1_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_12), .B1(f_s_Multiplier_0_1_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_4), .COUT(co_Multiplier_0_3_5), 
          .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1159[11] 1162[88])
    defparam Multiplier_0_add_3_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .B0(f_s_Multiplier_0_1_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_14), .B1(f_s_Multiplier_0_1_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_5), .COUT(co_Multiplier_0_3_6), 
          .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1168[11] 1171[88])
    defparam Multiplier_0_add_3_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .B0(f_s_Multiplier_0_1_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_16), .B1(f_s_Multiplier_0_1_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_6), .COUT(co_Multiplier_0_3_7), 
          .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1177[11] 1180[88])
    defparam Multiplier_0_add_3_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .B0(f_s_Multiplier_0_1_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(f_s_Multiplier_0_1_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_7), .COUT(co_Multiplier_0_3_8), 
          .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1186[11] 1189[88])
    defparam Multiplier_0_add_3_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_8.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_9 (.A0(GND_net), .B0(f_s_Multiplier_0_1_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(f_s_Multiplier_0_1_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
          .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1195[11] 1198[62])
    defparam Multiplier_0_add_3_9.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_9.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_9.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_9.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_10 (.A0(GND_net), .B0(f_s_Multiplier_0_1_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
          .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1204[11] 1207[63])
    defparam Multiplier_0_add_3_10.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_10.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_10.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_10.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_3_11 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1213[11] 1216[24])
    defparam Cadd_Multiplier_0_3_11.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_11.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_11.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_3_11.INJECT1_1 = "NO";
    CCU2C Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(s_Multiplier_0_3_8), .B1(f_Multiplier_0_pp_4_8), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_t_Multiplier_0_4_1), .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1222[11] 1224[100])
    defparam Cadd_t_Multiplier_0_4_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_t_Multiplier_0_4_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_t_Multiplier_0_4_1.INJECT1_0 = "NO";
    defparam Cadd_t_Multiplier_0_4_1.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .B0(f_Multiplier_0_pp_4_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_10), .B1(f_s_Multiplier_0_2_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_1), .COUT(co_t_Multiplier_0_4_2), 
          .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1230[11] 1233[69])
    defparam t_Multiplier_0_add_4_2.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_2.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_2.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_2.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .B0(f_s_Multiplier_0_2_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_12), .B1(f_s_Multiplier_0_2_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_2), .COUT(co_t_Multiplier_0_4_3), 
          .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1239[11] 1242[70])
    defparam t_Multiplier_0_add_4_3.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_3.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_3.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_3.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .B0(f_s_Multiplier_0_2_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_14), .B1(f_s_Multiplier_0_2_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_3), .COUT(co_t_Multiplier_0_4_4), 
          .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1248[11] 1251[70])
    defparam t_Multiplier_0_add_4_4.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_4.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_4.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_4.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .B0(f_s_Multiplier_0_2_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_16), .B1(f_s_Multiplier_0_2_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_4), .COUT(co_t_Multiplier_0_4_5), 
          .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1257[11] 1260[70])
    defparam t_Multiplier_0_add_4_5.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_5.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_5.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_5.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .B0(f_s_Multiplier_0_2_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_18), .B1(f_s_Multiplier_0_2_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_5), .COUT(co_t_Multiplier_0_4_6), 
          .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1266[11] 1269[70])
    defparam t_Multiplier_0_add_4_6.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_6.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_6.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_6.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .B0(f_s_Multiplier_0_2_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_20), .B1(f_s_Multiplier_0_2_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_6), .COUT(co_t_Multiplier_0_4_7), 
          .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1275[11] 1278[70])
    defparam t_Multiplier_0_add_4_7.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_7.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_7.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_7.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .B0(f_s_Multiplier_0_2_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_22), .B1(f_s_Multiplier_0_2_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_7), .COUT(co_t_Multiplier_0_4_8), 
          .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1284[11] 1287[70])
    defparam t_Multiplier_0_add_4_8.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_8.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_8.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_8.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .B0(f_s_Multiplier_0_2_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_t_Multiplier_0_4_8), .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1293[11] 1296[45])
    defparam t_Multiplier_0_add_4_9.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_9.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_9.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_9.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_0 (.A0(regb_b_0), .B0(regb_b_1), .C0(rega_a_1), 
          .D0(regb_b_0), .A1(rega_a_1), .B1(regb_b_1), .C1(rega_a_2), 
          .D1(regb_b_0), .CIN(Multiplier_0_cin_lr_0), .COUT(mco), .S0(Multiplier_0_pp_0_1), 
          .S1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1302[11] 1305[20])
    defparam Multiplier_0_mult_0_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_1 (.A0(rega_a_2), .B0(regb_b_1), .C0(rega_a_3), 
          .D0(regb_b_0), .A1(rega_a_3), .B1(regb_b_1), .C1(rega_a_4), 
          .D1(regb_b_0), .CIN(mco), .COUT(mco_1), .S0(Multiplier_0_pp_0_3), 
          .S1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1311[11] 1313[85])
    defparam Multiplier_0_mult_0_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_2 (.A0(rega_a_4), .B0(regb_b_1), .C0(rega_a_5), 
          .D0(regb_b_0), .A1(rega_a_5), .B1(regb_b_1), .C1(rega_a_6), 
          .D1(regb_b_0), .CIN(mco_1), .COUT(mco_2), .S0(Multiplier_0_pp_0_5), 
          .S1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1319[11] 1322[22])
    defparam Multiplier_0_mult_0_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_3 (.A0(rega_a_6), .B0(regb_b_1), .C0(rega_a_7), 
          .D0(regb_b_0), .A1(rega_a_7), .B1(regb_b_1), .C1(rega_a_8), 
          .D1(regb_b_0), .CIN(mco_2), .COUT(mco_3), .S0(Multiplier_0_pp_0_7), 
          .S1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1328[11] 1331[22])
    defparam Multiplier_0_mult_0_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_4 (.A0(rega_a_8), .B0(regb_b_1), .C0(rega_a_9), 
          .D0(regb_b_0), .A1(rega_a_9), .B1(regb_b_1), .C1(rega_a_10), 
          .D1(regb_b_0), .CIN(mco_3), .COUT(mco_4), .S0(Multiplier_0_pp_0_9), 
          .S1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1337[11] 1340[22])
    defparam Multiplier_0_mult_0_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_5 (.A0(rega_a_10), .B0(regb_b_1), .C0(Multiplier_0_mult_0_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_0_5_n1), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(mco_4), .COUT(mfco), .S0(Multiplier_0_pp_0_11), 
          .S1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1346[11] 1349[48])
    defparam Multiplier_0_mult_0_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_0 (.A0(regb_b_0), .B0(regb_b_3), .C0(rega_a_1), 
          .D0(regb_b_2), .A1(rega_a_1), .B1(regb_b_3), .C1(rega_a_2), 
          .D1(regb_b_2), .CIN(Multiplier_0_cin_lr_2), .COUT(mco_5), .S0(Multiplier_0_pp_1_3), 
          .S1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1355[11] 1358[22])
    defparam Multiplier_0_mult_2_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_1 (.A0(rega_a_2), .B0(regb_b_3), .C0(rega_a_3), 
          .D0(regb_b_2), .A1(rega_a_3), .B1(regb_b_3), .C1(rega_a_4), 
          .D1(regb_b_2), .CIN(mco_5), .COUT(mco_6), .S0(Multiplier_0_pp_1_5), 
          .S1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1364[11] 1367[22])
    defparam Multiplier_0_mult_2_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_2 (.A0(rega_a_4), .B0(regb_b_3), .C0(rega_a_5), 
          .D0(regb_b_2), .A1(rega_a_5), .B1(regb_b_3), .C1(rega_a_6), 
          .D1(regb_b_2), .CIN(mco_6), .COUT(mco_7), .S0(Multiplier_0_pp_1_7), 
          .S1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1373[11] 1376[22])
    defparam Multiplier_0_mult_2_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_3 (.A0(rega_a_6), .B0(regb_b_3), .C0(rega_a_7), 
          .D0(regb_b_2), .A1(rega_a_7), .B1(regb_b_3), .C1(rega_a_8), 
          .D1(regb_b_2), .CIN(mco_7), .COUT(mco_8), .S0(Multiplier_0_pp_1_9), 
          .S1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1382[11] 1385[22])
    defparam Multiplier_0_mult_2_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_4 (.A0(rega_a_8), .B0(regb_b_3), .C0(rega_a_9), 
          .D0(regb_b_2), .A1(rega_a_9), .B1(regb_b_3), .C1(rega_a_10), 
          .D1(regb_b_2), .CIN(mco_8), .COUT(mco_9), .S0(Multiplier_0_pp_1_11), 
          .S1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1391[11] 1394[22])
    defparam Multiplier_0_mult_2_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_5 (.A0(rega_a_10), .B0(regb_b_3), .C0(Multiplier_0_mult_2_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_2_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_2), .CIN(mco_9), .COUT(mfco_1), .S0(Multiplier_0_pp_1_13), 
          .S1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1400[11] 1403[50])
    defparam Multiplier_0_mult_2_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_0 (.A0(regb_b_0), .B0(regb_b_5), .C0(rega_a_1), 
          .D0(regb_b_4), .A1(rega_a_1), .B1(regb_b_5), .C1(rega_a_2), 
          .D1(regb_b_4), .CIN(Multiplier_0_cin_lr_4), .COUT(mco_10), .S0(Multiplier_0_pp_2_5), 
          .S1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1409[11] 1412[23])
    defparam Multiplier_0_mult_4_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_1 (.A0(rega_a_2), .B0(regb_b_5), .C0(rega_a_3), 
          .D0(regb_b_4), .A1(rega_a_3), .B1(regb_b_5), .C1(rega_a_4), 
          .D1(regb_b_4), .CIN(mco_10), .COUT(mco_11), .S0(Multiplier_0_pp_2_7), 
          .S1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1418[11] 1421[23])
    defparam Multiplier_0_mult_4_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_2 (.A0(rega_a_4), .B0(regb_b_5), .C0(rega_a_5), 
          .D0(regb_b_4), .A1(rega_a_5), .B1(regb_b_5), .C1(rega_a_6), 
          .D1(regb_b_4), .CIN(mco_11), .COUT(mco_12), .S0(Multiplier_0_pp_2_9), 
          .S1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1427[11] 1430[23])
    defparam Multiplier_0_mult_4_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_3 (.A0(rega_a_6), .B0(regb_b_5), .C0(rega_a_7), 
          .D0(regb_b_4), .A1(rega_a_7), .B1(regb_b_5), .C1(rega_a_8), 
          .D1(regb_b_4), .CIN(mco_12), .COUT(mco_13), .S0(Multiplier_0_pp_2_11), 
          .S1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1436[11] 1439[23])
    defparam Multiplier_0_mult_4_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_4 (.A0(rega_a_8), .B0(regb_b_5), .C0(rega_a_9), 
          .D0(regb_b_4), .A1(rega_a_9), .B1(regb_b_5), .C1(rega_a_10), 
          .D1(regb_b_4), .CIN(mco_13), .COUT(mco_14), .S0(Multiplier_0_pp_2_13), 
          .S1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1445[11] 1448[23])
    defparam Multiplier_0_mult_4_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_5 (.A0(rega_a_10), .B0(regb_b_5), .C0(Multiplier_0_mult_4_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_4_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_4), .CIN(mco_14), .COUT(mfco_2), .S0(Multiplier_0_pp_2_15), 
          .S1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1454[11] 1457[50])
    defparam Multiplier_0_mult_4_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_0 (.A0(regb_b_0), .B0(regb_b_7), .C0(rega_a_1), 
          .D0(regb_b_6), .A1(rega_a_1), .B1(regb_b_7), .C1(rega_a_2), 
          .D1(regb_b_6), .CIN(Multiplier_0_cin_lr_6), .COUT(mco_15), .S0(Multiplier_0_pp_3_7), 
          .S1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1463[11] 1466[23])
    defparam Multiplier_0_mult_6_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_1 (.A0(rega_a_2), .B0(regb_b_7), .C0(rega_a_3), 
          .D0(regb_b_6), .A1(rega_a_3), .B1(regb_b_7), .C1(rega_a_4), 
          .D1(regb_b_6), .CIN(mco_15), .COUT(mco_16), .S0(Multiplier_0_pp_3_9), 
          .S1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1472[11] 1475[23])
    defparam Multiplier_0_mult_6_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_2 (.A0(rega_a_4), .B0(regb_b_7), .C0(rega_a_5), 
          .D0(regb_b_6), .A1(rega_a_5), .B1(regb_b_7), .C1(rega_a_6), 
          .D1(regb_b_6), .CIN(mco_16), .COUT(mco_17), .S0(Multiplier_0_pp_3_11), 
          .S1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1481[11] 1484[23])
    defparam Multiplier_0_mult_6_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_3 (.A0(rega_a_6), .B0(regb_b_7), .C0(rega_a_7), 
          .D0(regb_b_6), .A1(rega_a_7), .B1(regb_b_7), .C1(rega_a_8), 
          .D1(regb_b_6), .CIN(mco_17), .COUT(mco_18), .S0(Multiplier_0_pp_3_13), 
          .S1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1490[11] 1493[23])
    defparam Multiplier_0_mult_6_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_4 (.A0(rega_a_8), .B0(regb_b_7), .C0(rega_a_9), 
          .D0(regb_b_6), .A1(rega_a_9), .B1(regb_b_7), .C1(rega_a_10), 
          .D1(regb_b_6), .CIN(mco_18), .COUT(mco_19), .S0(Multiplier_0_pp_3_15), 
          .S1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1499[11] 1502[23])
    defparam Multiplier_0_mult_6_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_5 (.A0(rega_a_10), .B0(regb_b_7), .C0(Multiplier_0_mult_6_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_6_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_6), .CIN(mco_19), .COUT(mfco_3), .S0(Multiplier_0_pp_3_17), 
          .S1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1508[11] 1511[50])
    defparam Multiplier_0_mult_6_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_0 (.A0(regb_b_0), .B0(regb_b_9), .C0(rega_a_1), 
          .D0(regb_b_8), .A1(rega_a_1), .B1(regb_b_9), .C1(rega_a_2), 
          .D1(regb_b_8), .CIN(Multiplier_0_cin_lr_8), .COUT(mco_20), .S0(Multiplier_0_pp_4_9), 
          .S1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1517[11] 1520[23])
    defparam Multiplier_0_mult_8_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_1 (.A0(rega_a_2), .B0(regb_b_9), .C0(rega_a_3), 
          .D0(regb_b_8), .A1(rega_a_3), .B1(regb_b_9), .C1(rega_a_4), 
          .D1(regb_b_8), .CIN(mco_20), .COUT(mco_21), .S0(Multiplier_0_pp_4_11), 
          .S1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1526[11] 1529[23])
    defparam Multiplier_0_mult_8_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_2 (.A0(rega_a_4), .B0(regb_b_9), .C0(rega_a_5), 
          .D0(regb_b_8), .A1(rega_a_5), .B1(regb_b_9), .C1(rega_a_6), 
          .D1(regb_b_8), .CIN(mco_21), .COUT(mco_22), .S0(Multiplier_0_pp_4_13), 
          .S1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1535[11] 1538[23])
    defparam Multiplier_0_mult_8_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_3 (.A0(rega_a_6), .B0(regb_b_9), .C0(rega_a_7), 
          .D0(regb_b_8), .A1(rega_a_7), .B1(regb_b_9), .C1(rega_a_8), 
          .D1(regb_b_8), .CIN(mco_22), .COUT(mco_23), .S0(Multiplier_0_pp_4_15), 
          .S1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1544[11] 1547[23])
    defparam Multiplier_0_mult_8_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_4 (.A0(rega_a_8), .B0(regb_b_9), .C0(rega_a_9), 
          .D0(regb_b_8), .A1(rega_a_9), .B1(regb_b_9), .C1(rega_a_10), 
          .D1(regb_b_8), .CIN(mco_23), .COUT(mco_24), .S0(Multiplier_0_pp_4_17), 
          .S1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1553[11] 1556[23])
    defparam Multiplier_0_mult_8_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_5 (.A0(rega_a_10), .B0(regb_b_9), .C0(Multiplier_0_mult_8_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_8_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_8), .CIN(mco_24), .COUT(mfco_4), .S0(Multiplier_0_pp_4_19), 
          .S1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1562[11] 1565[50])
    defparam Multiplier_0_mult_8_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .B0(VCC_net), 
          .C0(rega_a_1), .D0(regb_b_10), .A1(Multiplier_0_mult_10_0_n1), 
          .B1(VCC_net), .C1(rega_a_2), .D1(regb_b_10), .CIN(Multiplier_0_cin_lr_10), 
          .COUT(mco_25), .S0(Multiplier_0_pp_5_11), .S1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1571[11] 1574[50])
    defparam Multiplier_0_mult_10_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .B0(VCC_net), 
          .C0(rega_a_3), .D0(regb_b_10), .A1(Multiplier_0_mult_10_1_n1), 
          .B1(VCC_net), .C1(rega_a_4), .D1(regb_b_10), .CIN(mco_25), 
          .COUT(mco_26), .S0(Multiplier_0_pp_5_13), .S1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1580[11] 1583[23])
    defparam Multiplier_0_mult_10_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .B0(VCC_net), 
          .C0(rega_a_5), .D0(regb_b_10), .A1(Multiplier_0_mult_10_2_n1), 
          .B1(VCC_net), .C1(rega_a_6), .D1(regb_b_10), .CIN(mco_26), 
          .COUT(mco_27), .S0(Multiplier_0_pp_5_15), .S1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1589[11] 1592[23])
    defparam Multiplier_0_mult_10_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .B0(VCC_net), 
          .C0(rega_a_7), .D0(regb_b_10), .A1(Multiplier_0_mult_10_3_n1), 
          .B1(VCC_net), .C1(rega_a_8), .D1(regb_b_10), .CIN(mco_27), 
          .COUT(mco_28), .S0(Multiplier_0_pp_5_17), .S1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1598[11] 1601[23])
    defparam Multiplier_0_mult_10_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .B0(VCC_net), 
          .C0(rega_a_9), .D0(regb_b_10), .A1(Multiplier_0_mult_10_4_n1), 
          .B1(VCC_net), .C1(rega_a_10), .D1(regb_b_10), .CIN(mco_28), 
          .COUT(mco_29), .S0(Multiplier_0_pp_5_19), .S1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1607[11] 1610[23])
    defparam Multiplier_0_mult_10_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .B0(VCC_net), 
          .C0(Multiplier_0_mult_10_5_n2), .D0(VCC_net), .A1(rega_a_11), 
          .B1(regb_b_11), .C1(GND_net), .D1(regb_b_10), .CIN(mco_29), 
          .COUT(mfco_5), .S0(Multiplier_0_pp_5_21), .S1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1620[11] 1623[50])
    defparam Multiplier_0_mult_10_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_5.INJECT1_1 = "NO";
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(376[10:72])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(77[14] 83[27])
    
endmodule
//
// Verilog Description of module Multiplier_U0
//

module Multiplier_U0 (CIC1_out_clkSin, VCC_net, GND_net, MultDataB, 
            MultResult1) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/top.v(89[6:21])
    
    wire regb_b_1, Multiplier_0_mult_0_5_n1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, regb_b_3, Multiplier_0_mult_2_5_n1, Multiplier_0_pp_2_4, 
        regb_b_4, regb_b_5, Multiplier_0_mult_4_5_n1, Multiplier_0_pp_3_6, 
        regb_b_6, regb_b_7, Multiplier_0_mult_6_5_n1, Multiplier_0_pp_4_8, 
        regb_b_8, regb_b_9, Multiplier_0_mult_8_5_n1, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_10, 
        s_Multiplier_0_3_9, co_Multiplier_0_3_5, s_Multiplier_0_3_12, 
        s_Multiplier_0_3_11, co_Multiplier_0_3_6, s_Multiplier_0_3_14, 
        s_Multiplier_0_3_13, co_Multiplier_0_3_7, s_Multiplier_0_3_16, 
        s_Multiplier_0_3_15, co_Multiplier_0_3_8, s_Multiplier_0_3_18, 
        s_Multiplier_0_3_17, co_Multiplier_0_3_9, s_Multiplier_0_3_20, 
        s_Multiplier_0_3_19, co_Multiplier_0_3_10, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_21, s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, 
        co_t_Multiplier_0_4_2, co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, 
        co_t_Multiplier_0_4_5, co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, 
        co_t_Multiplier_0_4_8, mco, mco_1, mco_2, mco_3, mco_4, 
        Multiplier_0_mult_0_5_n2, mco_5, mco_6, mco_7, mco_8, mco_9, 
        Multiplier_0_mult_2_5_n2, mco_10, mco_11, mco_12, mco_13, 
        mco_14, Multiplier_0_mult_4_5_n2, mco_15, mco_16, mco_17, 
        mco_18, mco_19, Multiplier_0_mult_6_5_n2, mco_20, mco_21, 
        mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, Multiplier_0_mult_10_0_n1, 
        mco_25, mco_26, mco_27, mco_28, mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    FD1P3DX FF_98 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataB[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    CCU2C Multiplier_0_cin_lr_add_0 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(788[11] 790[76])
    defparam Multiplier_0_cin_lr_add_0.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_0.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_0.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_0_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(796[11] 798[79])
    defparam Multiplier_0_Cadd_0_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_0_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_0_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_0_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_2 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(804[11] 806[76])
    defparam Multiplier_0_cin_lr_add_2.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_2.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_2.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_2_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(812[11] 815[17])
    defparam Multiplier_0_Cadd_2_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_2_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_2_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_2_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_4 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(821[11] 823[76])
    defparam Multiplier_0_cin_lr_add_4.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_4.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_4.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_4_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(829[11] 832[17])
    defparam Multiplier_0_Cadd_4_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_4_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_4_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_4_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_6 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(838[11] 840[76])
    defparam Multiplier_0_cin_lr_add_6.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_6.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_6.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_6_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(846[11] 849[17])
    defparam Multiplier_0_Cadd_6_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_6_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_6_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_6_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_8 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(855[11] 857[76])
    defparam Multiplier_0_cin_lr_add_8.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_8.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_8.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_8.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_8_6 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(863[11] 866[17])
    defparam Multiplier_0_Cadd_8_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_8_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_8_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_8_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_cin_lr_add_10 (.A0(VCC_net), .B0(VCC_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), 
          .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(872[11] 874[77])
    defparam Multiplier_0_cin_lr_add_10.INIT0 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_10.INIT1 = 16'b0000000000000000;
    defparam Multiplier_0_cin_lr_add_10.INJECT1_0 = "NO";
    defparam Multiplier_0_cin_lr_add_10.INJECT1_1 = "NO";
    CCU2C Multiplier_0_Cadd_10_6 (.A0(VCC_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(880[11] 883[17])
    defparam Multiplier_0_Cadd_10_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_10_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_Cadd_10_6.INJECT1_0 = "NO";
    defparam Multiplier_0_Cadd_10_6.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_0_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(Multiplier_0_pp_0_2), .B1(Multiplier_0_pp_1_2), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_0_1), .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(889[11] 892[36])
    defparam Cadd_Multiplier_0_0_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_0_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .B0(Multiplier_0_pp_1_3), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_4), .B1(Multiplier_0_pp_1_4), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_1), .COUT(co_Multiplier_0_0_2), 
          .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(898[11] 901[86])
    defparam Multiplier_0_add_0_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .B0(Multiplier_0_pp_1_5), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_6), .B1(Multiplier_0_pp_1_6), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_2), .COUT(co_Multiplier_0_0_3), 
          .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(907[11] 910[86])
    defparam Multiplier_0_add_0_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .B0(Multiplier_0_pp_1_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_8), .B1(Multiplier_0_pp_1_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_3), .COUT(co_Multiplier_0_0_4), 
          .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(916[11] 919[86])
    defparam Multiplier_0_add_0_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .B0(Multiplier_0_pp_1_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_10), .B1(Multiplier_0_pp_1_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_4), .COUT(co_Multiplier_0_0_5), 
          .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(925[11] 928[87])
    defparam Multiplier_0_add_0_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .B0(Multiplier_0_pp_1_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_0_12), .B1(Multiplier_0_pp_1_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_5), .COUT(co_Multiplier_0_0_6), 
          .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(934[11] 937[88])
    defparam Multiplier_0_add_0_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .B0(Multiplier_0_pp_1_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(Multiplier_0_pp_1_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_0_6), .COUT(co_Multiplier_0_0_7), 
          .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(943[11] 946[88])
    defparam Multiplier_0_add_0_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_0_8 (.A0(GND_net), .B0(Multiplier_0_pp_1_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
          .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(952[11] 955[62])
    defparam Multiplier_0_add_0_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_0_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_0_8.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_0_9 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(961[11] 964[24])
    defparam Cadd_Multiplier_0_0_9.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_9.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_0_9.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_0_9.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_1_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(Multiplier_0_pp_2_6), .B1(Multiplier_0_pp_3_6), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_1_1), .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(970[11] 973[36])
    defparam Cadd_Multiplier_0_1_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_1_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .B0(Multiplier_0_pp_3_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_8), .B1(Multiplier_0_pp_3_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_1), .COUT(co_Multiplier_0_1_2), 
          .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(979[11] 982[86])
    defparam Multiplier_0_add_1_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .B0(Multiplier_0_pp_3_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_10), .B1(Multiplier_0_pp_3_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_2), .COUT(co_Multiplier_0_1_3), 
          .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(988[11] 991[87])
    defparam Multiplier_0_add_1_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .B0(Multiplier_0_pp_3_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_12), .B1(Multiplier_0_pp_3_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_3), .COUT(co_Multiplier_0_1_4), 
          .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(997[11] 1000[88])
    defparam Multiplier_0_add_1_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .B0(Multiplier_0_pp_3_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_14), .B1(Multiplier_0_pp_3_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_4), .COUT(co_Multiplier_0_1_5), 
          .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1006[11] 1009[88])
    defparam Multiplier_0_add_1_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .B0(Multiplier_0_pp_3_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_2_16), .B1(Multiplier_0_pp_3_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_5), .COUT(co_Multiplier_0_1_6), 
          .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1015[11] 1018[88])
    defparam Multiplier_0_add_1_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .B0(Multiplier_0_pp_3_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(Multiplier_0_pp_3_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_1_6), .COUT(co_Multiplier_0_1_7), 
          .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1024[11] 1027[88])
    defparam Multiplier_0_add_1_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_1_8 (.A0(GND_net), .B0(Multiplier_0_pp_3_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
          .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1033[11] 1036[62])
    defparam Multiplier_0_add_1_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_1_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_1_8.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_1_9 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1042[11] 1045[24])
    defparam Cadd_Multiplier_0_1_9.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_9.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_1_9.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_1_9.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_2_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(Multiplier_0_pp_4_10), .B1(Multiplier_0_pp_5_10), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_2_1), .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1051[11] 1054[36])
    defparam Cadd_Multiplier_0_2_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_2_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_2_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_2_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .B0(Multiplier_0_pp_5_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_12), .B1(Multiplier_0_pp_5_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_1), .COUT(co_Multiplier_0_2_2), 
          .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1060[11] 1063[88])
    defparam Multiplier_0_add_2_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .B0(Multiplier_0_pp_5_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_14), .B1(Multiplier_0_pp_5_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_2), .COUT(co_Multiplier_0_2_3), 
          .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1069[11] 1072[88])
    defparam Multiplier_0_add_2_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .B0(Multiplier_0_pp_5_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_16), .B1(Multiplier_0_pp_5_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_3), .COUT(co_Multiplier_0_2_4), 
          .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1078[11] 1081[88])
    defparam Multiplier_0_add_2_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .B0(Multiplier_0_pp_5_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_18), .B1(Multiplier_0_pp_5_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_4), .COUT(co_Multiplier_0_2_5), 
          .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1087[11] 1090[88])
    defparam Multiplier_0_add_2_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .B0(Multiplier_0_pp_5_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(Multiplier_0_pp_4_20), .B1(Multiplier_0_pp_5_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_5), .COUT(co_Multiplier_0_2_6), 
          .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1096[11] 1099[88])
    defparam Multiplier_0_add_2_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .B0(Multiplier_0_pp_5_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(Multiplier_0_pp_5_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_2_6), .COUT(co_Multiplier_0_2_7), 
          .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1105[11] 1108[88])
    defparam Multiplier_0_add_2_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_2_8 (.A0(GND_net), .B0(Multiplier_0_pp_5_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1114[11] 1117[43])
    defparam Multiplier_0_add_2_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_2_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_2_8.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_3_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(f_s_Multiplier_0_0_4), .B1(f_Multiplier_0_pp_2_4), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_Multiplier_0_3_1), .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1123[11] 1126[36])
    defparam Cadd_Multiplier_0_3_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_1.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_3_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .B0(f_Multiplier_0_pp_2_5), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_6), .B1(f_s_Multiplier_0_1_6), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_1), .COUT(co_Multiplier_0_3_2), 
          .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1132[11] 1135[86])
    defparam Multiplier_0_add_3_2.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_2.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_2.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .B0(f_s_Multiplier_0_1_7), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_8), .B1(f_s_Multiplier_0_1_8), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_2), .COUT(co_Multiplier_0_3_3), 
          .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1141[11] 1144[86])
    defparam Multiplier_0_add_3_3.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_3.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_3.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .B0(f_s_Multiplier_0_1_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_10), .B1(f_s_Multiplier_0_1_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_3), .COUT(co_Multiplier_0_3_4), 
          .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1150[11] 1153[87])
    defparam Multiplier_0_add_3_4.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_4.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_4.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .B0(f_s_Multiplier_0_1_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_12), .B1(f_s_Multiplier_0_1_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_4), .COUT(co_Multiplier_0_3_5), 
          .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1159[11] 1162[88])
    defparam Multiplier_0_add_3_5.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_5.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_5.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .B0(f_s_Multiplier_0_1_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_14), .B1(f_s_Multiplier_0_1_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_5), .COUT(co_Multiplier_0_3_6), 
          .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1168[11] 1171[88])
    defparam Multiplier_0_add_3_6.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_6.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_6.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_6.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .B0(f_s_Multiplier_0_1_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(f_s_Multiplier_0_0_16), .B1(f_s_Multiplier_0_1_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_6), .COUT(co_Multiplier_0_3_7), 
          .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1177[11] 1180[88])
    defparam Multiplier_0_add_3_7.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_7.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_7.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_7.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .B0(f_s_Multiplier_0_1_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(f_s_Multiplier_0_1_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_7), .COUT(co_Multiplier_0_3_8), 
          .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1186[11] 1189[88])
    defparam Multiplier_0_add_3_8.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_8.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_8.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_8.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_9 (.A0(GND_net), .B0(f_s_Multiplier_0_1_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(f_s_Multiplier_0_1_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
          .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1195[11] 1198[62])
    defparam Multiplier_0_add_3_9.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_9.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_9.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_9.INJECT1_1 = "NO";
    CCU2C Multiplier_0_add_3_10 (.A0(GND_net), .B0(f_s_Multiplier_0_1_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
          .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1204[11] 1207[63])
    defparam Multiplier_0_add_3_10.INIT0 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_10.INIT1 = 16'b0110011010101010;
    defparam Multiplier_0_add_3_10.INJECT1_0 = "NO";
    defparam Multiplier_0_add_3_10.INJECT1_1 = "NO";
    CCU2C Cadd_Multiplier_0_3_11 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1213[11] 1216[24])
    defparam Cadd_Multiplier_0_3_11.INIT0 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_11.INIT1 = 16'b0110011010101010;
    defparam Cadd_Multiplier_0_3_11.INJECT1_0 = "NO";
    defparam Cadd_Multiplier_0_3_11.INJECT1_1 = "NO";
    CCU2C Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(s_Multiplier_0_3_8), .B1(f_Multiplier_0_pp_4_8), 
          .C1(VCC_net), .D1(VCC_net), .COUT(co_t_Multiplier_0_4_1), .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1222[11] 1224[100])
    defparam Cadd_t_Multiplier_0_4_1.INIT0 = 16'b0110011010101010;
    defparam Cadd_t_Multiplier_0_4_1.INIT1 = 16'b0110011010101010;
    defparam Cadd_t_Multiplier_0_4_1.INJECT1_0 = "NO";
    defparam Cadd_t_Multiplier_0_4_1.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .B0(f_Multiplier_0_pp_4_9), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_10), .B1(f_s_Multiplier_0_2_10), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_1), .COUT(co_t_Multiplier_0_4_2), 
          .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1230[11] 1233[69])
    defparam t_Multiplier_0_add_4_2.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_2.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_2.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_2.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .B0(f_s_Multiplier_0_2_11), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_12), .B1(f_s_Multiplier_0_2_12), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_2), .COUT(co_t_Multiplier_0_4_3), 
          .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1239[11] 1242[70])
    defparam t_Multiplier_0_add_4_3.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_3.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_3.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_3.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .B0(f_s_Multiplier_0_2_13), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_14), .B1(f_s_Multiplier_0_2_14), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_3), .COUT(co_t_Multiplier_0_4_4), 
          .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1248[11] 1251[70])
    defparam t_Multiplier_0_add_4_4.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_4.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_4.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_4.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .B0(f_s_Multiplier_0_2_15), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_16), .B1(f_s_Multiplier_0_2_16), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_4), .COUT(co_t_Multiplier_0_4_5), 
          .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1257[11] 1260[70])
    defparam t_Multiplier_0_add_4_5.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_5.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_5.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_5.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .B0(f_s_Multiplier_0_2_17), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_18), .B1(f_s_Multiplier_0_2_18), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_5), .COUT(co_t_Multiplier_0_4_6), 
          .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1266[11] 1269[70])
    defparam t_Multiplier_0_add_4_6.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_6.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_6.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_6.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .B0(f_s_Multiplier_0_2_19), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_20), .B1(f_s_Multiplier_0_2_20), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_6), .COUT(co_t_Multiplier_0_4_7), 
          .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1275[11] 1278[70])
    defparam t_Multiplier_0_add_4_7.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_7.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_7.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_7.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .B0(f_s_Multiplier_0_2_21), 
          .C0(VCC_net), .D0(VCC_net), .A1(s_Multiplier_0_3_22), .B1(f_s_Multiplier_0_2_22), 
          .C1(VCC_net), .D1(VCC_net), .CIN(co_t_Multiplier_0_4_7), .COUT(co_t_Multiplier_0_4_8), 
          .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1284[11] 1287[70])
    defparam t_Multiplier_0_add_4_8.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_8.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_8.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_8.INJECT1_1 = "NO";
    CCU2C t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .B0(f_s_Multiplier_0_2_23), 
          .C0(VCC_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co_t_Multiplier_0_4_8), .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1293[11] 1296[45])
    defparam t_Multiplier_0_add_4_9.INIT0 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_9.INIT1 = 16'b0110011010101010;
    defparam t_Multiplier_0_add_4_9.INJECT1_0 = "NO";
    defparam t_Multiplier_0_add_4_9.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_0 (.A0(regb_b_0), .B0(regb_b_1), .C0(rega_a_1), 
          .D0(regb_b_0), .A1(rega_a_1), .B1(regb_b_1), .C1(rega_a_2), 
          .D1(regb_b_0), .CIN(Multiplier_0_cin_lr_0), .COUT(mco), .S0(Multiplier_0_pp_0_1), 
          .S1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1302[11] 1305[20])
    defparam Multiplier_0_mult_0_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_1 (.A0(rega_a_2), .B0(regb_b_1), .C0(rega_a_3), 
          .D0(regb_b_0), .A1(rega_a_3), .B1(regb_b_1), .C1(rega_a_4), 
          .D1(regb_b_0), .CIN(mco), .COUT(mco_1), .S0(Multiplier_0_pp_0_3), 
          .S1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1311[11] 1313[85])
    defparam Multiplier_0_mult_0_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_2 (.A0(rega_a_4), .B0(regb_b_1), .C0(rega_a_5), 
          .D0(regb_b_0), .A1(rega_a_5), .B1(regb_b_1), .C1(rega_a_6), 
          .D1(regb_b_0), .CIN(mco_1), .COUT(mco_2), .S0(Multiplier_0_pp_0_5), 
          .S1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1319[11] 1322[22])
    defparam Multiplier_0_mult_0_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_3 (.A0(rega_a_6), .B0(regb_b_1), .C0(rega_a_7), 
          .D0(regb_b_0), .A1(rega_a_7), .B1(regb_b_1), .C1(rega_a_8), 
          .D1(regb_b_0), .CIN(mco_2), .COUT(mco_3), .S0(Multiplier_0_pp_0_7), 
          .S1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1328[11] 1331[22])
    defparam Multiplier_0_mult_0_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_4 (.A0(rega_a_8), .B0(regb_b_1), .C0(rega_a_9), 
          .D0(regb_b_0), .A1(rega_a_9), .B1(regb_b_1), .C1(rega_a_10), 
          .D1(regb_b_0), .CIN(mco_3), .COUT(mco_4), .S0(Multiplier_0_pp_0_9), 
          .S1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1337[11] 1340[22])
    defparam Multiplier_0_mult_0_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_0_5 (.A0(rega_a_10), .B0(regb_b_1), .C0(Multiplier_0_mult_0_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_0_5_n1), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(mco_4), .COUT(mfco), .S0(Multiplier_0_pp_0_11), 
          .S1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1346[11] 1349[48])
    defparam Multiplier_0_mult_0_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_0_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_0_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_0 (.A0(regb_b_0), .B0(regb_b_3), .C0(rega_a_1), 
          .D0(regb_b_2), .A1(rega_a_1), .B1(regb_b_3), .C1(rega_a_2), 
          .D1(regb_b_2), .CIN(Multiplier_0_cin_lr_2), .COUT(mco_5), .S0(Multiplier_0_pp_1_3), 
          .S1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1355[11] 1358[22])
    defparam Multiplier_0_mult_2_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_1 (.A0(rega_a_2), .B0(regb_b_3), .C0(rega_a_3), 
          .D0(regb_b_2), .A1(rega_a_3), .B1(regb_b_3), .C1(rega_a_4), 
          .D1(regb_b_2), .CIN(mco_5), .COUT(mco_6), .S0(Multiplier_0_pp_1_5), 
          .S1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1364[11] 1367[22])
    defparam Multiplier_0_mult_2_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_2 (.A0(rega_a_4), .B0(regb_b_3), .C0(rega_a_5), 
          .D0(regb_b_2), .A1(rega_a_5), .B1(regb_b_3), .C1(rega_a_6), 
          .D1(regb_b_2), .CIN(mco_6), .COUT(mco_7), .S0(Multiplier_0_pp_1_7), 
          .S1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1373[11] 1376[22])
    defparam Multiplier_0_mult_2_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_3 (.A0(rega_a_6), .B0(regb_b_3), .C0(rega_a_7), 
          .D0(regb_b_2), .A1(rega_a_7), .B1(regb_b_3), .C1(rega_a_8), 
          .D1(regb_b_2), .CIN(mco_7), .COUT(mco_8), .S0(Multiplier_0_pp_1_9), 
          .S1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1382[11] 1385[22])
    defparam Multiplier_0_mult_2_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_4 (.A0(rega_a_8), .B0(regb_b_3), .C0(rega_a_9), 
          .D0(regb_b_2), .A1(rega_a_9), .B1(regb_b_3), .C1(rega_a_10), 
          .D1(regb_b_2), .CIN(mco_8), .COUT(mco_9), .S0(Multiplier_0_pp_1_11), 
          .S1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1391[11] 1394[22])
    defparam Multiplier_0_mult_2_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_2_5 (.A0(rega_a_10), .B0(regb_b_3), .C0(Multiplier_0_mult_2_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_2_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_2), .CIN(mco_9), .COUT(mfco_1), .S0(Multiplier_0_pp_1_13), 
          .S1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1400[11] 1403[50])
    defparam Multiplier_0_mult_2_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_2_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_2_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_0 (.A0(regb_b_0), .B0(regb_b_5), .C0(rega_a_1), 
          .D0(regb_b_4), .A1(rega_a_1), .B1(regb_b_5), .C1(rega_a_2), 
          .D1(regb_b_4), .CIN(Multiplier_0_cin_lr_4), .COUT(mco_10), .S0(Multiplier_0_pp_2_5), 
          .S1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1409[11] 1412[23])
    defparam Multiplier_0_mult_4_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_1 (.A0(rega_a_2), .B0(regb_b_5), .C0(rega_a_3), 
          .D0(regb_b_4), .A1(rega_a_3), .B1(regb_b_5), .C1(rega_a_4), 
          .D1(regb_b_4), .CIN(mco_10), .COUT(mco_11), .S0(Multiplier_0_pp_2_7), 
          .S1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1418[11] 1421[23])
    defparam Multiplier_0_mult_4_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_2 (.A0(rega_a_4), .B0(regb_b_5), .C0(rega_a_5), 
          .D0(regb_b_4), .A1(rega_a_5), .B1(regb_b_5), .C1(rega_a_6), 
          .D1(regb_b_4), .CIN(mco_11), .COUT(mco_12), .S0(Multiplier_0_pp_2_9), 
          .S1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1427[11] 1430[23])
    defparam Multiplier_0_mult_4_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_3 (.A0(rega_a_6), .B0(regb_b_5), .C0(rega_a_7), 
          .D0(regb_b_4), .A1(rega_a_7), .B1(regb_b_5), .C1(rega_a_8), 
          .D1(regb_b_4), .CIN(mco_12), .COUT(mco_13), .S0(Multiplier_0_pp_2_11), 
          .S1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1436[11] 1439[23])
    defparam Multiplier_0_mult_4_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_4 (.A0(rega_a_8), .B0(regb_b_5), .C0(rega_a_9), 
          .D0(regb_b_4), .A1(rega_a_9), .B1(regb_b_5), .C1(rega_a_10), 
          .D1(regb_b_4), .CIN(mco_13), .COUT(mco_14), .S0(Multiplier_0_pp_2_13), 
          .S1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1445[11] 1448[23])
    defparam Multiplier_0_mult_4_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_4_5 (.A0(rega_a_10), .B0(regb_b_5), .C0(Multiplier_0_mult_4_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_4_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_4), .CIN(mco_14), .COUT(mfco_2), .S0(Multiplier_0_pp_2_15), 
          .S1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1454[11] 1457[50])
    defparam Multiplier_0_mult_4_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_4_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_4_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_0 (.A0(regb_b_0), .B0(regb_b_7), .C0(rega_a_1), 
          .D0(regb_b_6), .A1(rega_a_1), .B1(regb_b_7), .C1(rega_a_2), 
          .D1(regb_b_6), .CIN(Multiplier_0_cin_lr_6), .COUT(mco_15), .S0(Multiplier_0_pp_3_7), 
          .S1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1463[11] 1466[23])
    defparam Multiplier_0_mult_6_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_1 (.A0(rega_a_2), .B0(regb_b_7), .C0(rega_a_3), 
          .D0(regb_b_6), .A1(rega_a_3), .B1(regb_b_7), .C1(rega_a_4), 
          .D1(regb_b_6), .CIN(mco_15), .COUT(mco_16), .S0(Multiplier_0_pp_3_9), 
          .S1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1472[11] 1475[23])
    defparam Multiplier_0_mult_6_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_2 (.A0(rega_a_4), .B0(regb_b_7), .C0(rega_a_5), 
          .D0(regb_b_6), .A1(rega_a_5), .B1(regb_b_7), .C1(rega_a_6), 
          .D1(regb_b_6), .CIN(mco_16), .COUT(mco_17), .S0(Multiplier_0_pp_3_11), 
          .S1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1481[11] 1484[23])
    defparam Multiplier_0_mult_6_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_3 (.A0(rega_a_6), .B0(regb_b_7), .C0(rega_a_7), 
          .D0(regb_b_6), .A1(rega_a_7), .B1(regb_b_7), .C1(rega_a_8), 
          .D1(regb_b_6), .CIN(mco_17), .COUT(mco_18), .S0(Multiplier_0_pp_3_13), 
          .S1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1490[11] 1493[23])
    defparam Multiplier_0_mult_6_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_4 (.A0(rega_a_8), .B0(regb_b_7), .C0(rega_a_9), 
          .D0(regb_b_6), .A1(rega_a_9), .B1(regb_b_7), .C1(rega_a_10), 
          .D1(regb_b_6), .CIN(mco_18), .COUT(mco_19), .S0(Multiplier_0_pp_3_15), 
          .S1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1499[11] 1502[23])
    defparam Multiplier_0_mult_6_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_6_5 (.A0(rega_a_10), .B0(regb_b_7), .C0(Multiplier_0_mult_6_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_6_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_6), .CIN(mco_19), .COUT(mfco_3), .S0(Multiplier_0_pp_3_17), 
          .S1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1508[11] 1511[50])
    defparam Multiplier_0_mult_6_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_6_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_6_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_0 (.A0(regb_b_0), .B0(regb_b_9), .C0(rega_a_1), 
          .D0(regb_b_8), .A1(rega_a_1), .B1(regb_b_9), .C1(rega_a_2), 
          .D1(regb_b_8), .CIN(Multiplier_0_cin_lr_8), .COUT(mco_20), .S0(Multiplier_0_pp_4_9), 
          .S1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1517[11] 1520[23])
    defparam Multiplier_0_mult_8_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_1 (.A0(rega_a_2), .B0(regb_b_9), .C0(rega_a_3), 
          .D0(regb_b_8), .A1(rega_a_3), .B1(regb_b_9), .C1(rega_a_4), 
          .D1(regb_b_8), .CIN(mco_20), .COUT(mco_21), .S0(Multiplier_0_pp_4_11), 
          .S1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1526[11] 1529[23])
    defparam Multiplier_0_mult_8_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_2 (.A0(rega_a_4), .B0(regb_b_9), .C0(rega_a_5), 
          .D0(regb_b_8), .A1(rega_a_5), .B1(regb_b_9), .C1(rega_a_6), 
          .D1(regb_b_8), .CIN(mco_21), .COUT(mco_22), .S0(Multiplier_0_pp_4_13), 
          .S1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1535[11] 1538[23])
    defparam Multiplier_0_mult_8_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_3 (.A0(rega_a_6), .B0(regb_b_9), .C0(rega_a_7), 
          .D0(regb_b_8), .A1(rega_a_7), .B1(regb_b_9), .C1(rega_a_8), 
          .D1(regb_b_8), .CIN(mco_22), .COUT(mco_23), .S0(Multiplier_0_pp_4_15), 
          .S1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1544[11] 1547[23])
    defparam Multiplier_0_mult_8_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_4 (.A0(rega_a_8), .B0(regb_b_9), .C0(rega_a_9), 
          .D0(regb_b_8), .A1(rega_a_9), .B1(regb_b_9), .C1(rega_a_10), 
          .D1(regb_b_8), .CIN(mco_23), .COUT(mco_24), .S0(Multiplier_0_pp_4_17), 
          .S1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1553[11] 1556[23])
    defparam Multiplier_0_mult_8_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_8_5 (.A0(rega_a_10), .B0(regb_b_9), .C0(Multiplier_0_mult_8_5_n2), 
          .D0(VCC_net), .A1(Multiplier_0_mult_8_5_n1), .B1(VCC_net), .C1(GND_net), 
          .D1(regb_b_8), .CIN(mco_24), .COUT(mfco_4), .S0(Multiplier_0_pp_4_19), 
          .S1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1562[11] 1565[50])
    defparam Multiplier_0_mult_8_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_8_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_8_5.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .B0(VCC_net), 
          .C0(rega_a_1), .D0(regb_b_10), .A1(Multiplier_0_mult_10_0_n1), 
          .B1(VCC_net), .C1(rega_a_2), .D1(regb_b_10), .CIN(Multiplier_0_cin_lr_10), 
          .COUT(mco_25), .S0(Multiplier_0_pp_5_11), .S1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1571[11] 1574[50])
    defparam Multiplier_0_mult_10_0.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_0.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_0.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_0.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .B0(VCC_net), 
          .C0(rega_a_3), .D0(regb_b_10), .A1(Multiplier_0_mult_10_1_n1), 
          .B1(VCC_net), .C1(rega_a_4), .D1(regb_b_10), .CIN(mco_25), 
          .COUT(mco_26), .S0(Multiplier_0_pp_5_13), .S1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1580[11] 1583[23])
    defparam Multiplier_0_mult_10_1.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_1.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_1.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_1.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .B0(VCC_net), 
          .C0(rega_a_5), .D0(regb_b_10), .A1(Multiplier_0_mult_10_2_n1), 
          .B1(VCC_net), .C1(rega_a_6), .D1(regb_b_10), .CIN(mco_26), 
          .COUT(mco_27), .S0(Multiplier_0_pp_5_15), .S1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1589[11] 1592[23])
    defparam Multiplier_0_mult_10_2.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_2.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_2.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_2.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .B0(VCC_net), 
          .C0(rega_a_7), .D0(regb_b_10), .A1(Multiplier_0_mult_10_3_n1), 
          .B1(VCC_net), .C1(rega_a_8), .D1(regb_b_10), .CIN(mco_27), 
          .COUT(mco_28), .S0(Multiplier_0_pp_5_17), .S1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1598[11] 1601[23])
    defparam Multiplier_0_mult_10_3.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_3.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_3.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_3.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .B0(VCC_net), 
          .C0(rega_a_9), .D0(regb_b_10), .A1(Multiplier_0_mult_10_4_n1), 
          .B1(VCC_net), .C1(rega_a_10), .D1(regb_b_10), .CIN(mco_28), 
          .COUT(mco_29), .S0(Multiplier_0_pp_5_19), .S1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1607[11] 1610[23])
    defparam Multiplier_0_mult_10_4.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_4.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_4.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_4.INJECT1_1 = "NO";
    CCU2C Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .B0(VCC_net), 
          .C0(Multiplier_0_mult_10_5_n2), .D0(VCC_net), .A1(rega_a_11), 
          .B1(regb_b_11), .C1(GND_net), .D1(regb_b_10), .CIN(mco_29), 
          .COUT(mfco_5), .S0(Multiplier_0_pp_5_21), .S1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(1620[11] 1623[50])
    defparam Multiplier_0_mult_10_5.INIT0 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_5.INIT1 = 16'b0111100010001000;
    defparam Multiplier_0_mult_10_5.INJECT1_0 = "NO";
    defparam Multiplier_0_mult_10_5.INJECT1_1 = "NO";
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/IP/Multiplier/Multiplier.v(376[10:72])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/Master Thesis/1bitSDR/1bitSDRLatticeTest/First_Implementation/source/AMDemod.v(69[14] 75[27])
    
endmodule
