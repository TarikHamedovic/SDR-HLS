// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Thu Oct 31 10:30:10 2024
//
// Verilog Description of module top
//

module top (osc_clk, i_Rx_Serial, o_Tx_Serial, MYLED, XOut, RFIn, 
            DiffOut, PWMOut, PWMOutP1, PWMOutP2, PWMOutP3, PWMOutP4, 
            PWMOutN1, PWMOutN2, PWMOutN3, PWMOutN4, sinGen, sin_out, 
            CIC_out_clkSin) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(45[8:11])
    input osc_clk;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(47[13:20])
    input i_Rx_Serial;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(48[13:24])
    output o_Tx_Serial;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(49[11:22])
    output [7:0]MYLED;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    output XOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(54[9:13])
    input RFIn;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(55[9:13])
    output DiffOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(56[9:16])
    output PWMOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(57[9:15])
    output PWMOutP1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(58[9:17])
    output PWMOutP2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(59[9:17])
    output PWMOutP3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(60[9:17])
    output PWMOutP4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(61[9:17])
    output PWMOutN1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(62[9:17])
    output PWMOutN2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(63[9:17])
    output PWMOutN3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(64[9:17])
    output PWMOutN4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(65[9:17])
    output sinGen;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(66[9:15])
    output sin_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(67[9:16])
    output CIC_out_clkSin;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(68[9:23])
    
    wire osc_clk_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(47[13:20])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(86[6:21])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, MYLED_0_6, MYLED_0_5, MYLED_0_4, 
        MYLED_0_3, MYLED_0_2, MYLED_0_1, MYLED_0_0, RFIn_c, DiffOut_c, 
        PWMOutP4_c, PWMOutN4_c, sinGen_c, o_Rx_DV;
    wire [7:0]o_Rx_Byte;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(74[10:19])
    
    wire o_Rx_DV1;
    wire [7:0]o_Rx_Byte1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(77[11:21])
    wire [11:0]MixerOutSin;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(82[20:31])
    wire [11:0]MixerOutCos;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(83[20:31])
    wire [11:0]CIC1_outSin;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(85[20:31])
    wire [11:0]CIC1_outCos;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(88[20:31])
    wire [63:0]phase_accum;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(90[13:24])
    wire [12:0]LOSine;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(91[20:26])
    wire [12:0]LOCosine;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(92[20:28])
    wire [63:0]phase_inc_carrGen;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(94[19:36])
    wire [63:0]phase_inc_carrGen1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(95[19:37])
    wire [11:0]DemodOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(98[20:28])
    
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire [7:0]CICGain;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(100[11:18])
    
    wire n16276, n180, n7, n6, n5, n4, n3, n2, n37, n36, 
        n35, n34, n33, n32_adj_2749, n31_adj_2750, n30_adj_2751, 
        n29_adj_2752, n28_adj_2753, n27_adj_2754, n26_adj_2755, n25_adj_2756, 
        n24, n23, n22, n21, n20, n19, n18, n17, n2563, n16058, 
        n2331, n16, n15, n14, n13, n12, n11, n10, n9, n8, 
        n7_adj_2757, n6_adj_2758, n5_adj_2759, n4_adj_2760, n3_adj_2761, 
        n2_adj_2762, n16275, n177, n16056, n16055, n16274, n16273, 
        n16272, n16266, n16265, n16264, n16263, n16262, n16261, 
        n16260, n16259, n16258, n16252, n16251, n16250, n16249, 
        n16248, n16247, n16246, n16245, n2392, n16244, n2387, 
        n16238, n16237, n16236, n16235, n2381, n16234, n16233, 
        n16232, n16231, n16230, n15839, cout;
    wire [63:0]phase_accum_adj_5658;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(29[19:30])
    
    wire n90, n87, n84, n81, n78;
    wire [11:0]MixerOutSin_11__N_236;
    wire [11:0]MixerOutCos_11__N_250;
    
    wire n174;
    wire [71:0]d_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(30[26:31])
    wire [71:0]d_d_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(30[33:40])
    wire [71:0]d1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(35[26:28])
    wire [71:0]d2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(36[26:28])
    wire [71:0]d3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(37[26:28])
    wire [71:0]d4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(38[26:28])
    wire [71:0]d5;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(39[26:28])
    wire [71:0]d6;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(43[26:28])
    wire [71:0]d_d6;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(43[30:34])
    wire [71:0]d7;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(44[26:28])
    wire [71:0]d_d7;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(44[30:34])
    wire [71:0]d8;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(45[26:28])
    wire [71:0]d_d8;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(45[30:34])
    wire [71:0]d9;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(46[26:28])
    wire [71:0]d_d9;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(46[30:34])
    
    wire n16054, n171, n15913;
    wire [15:0]count;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(50[14:19])
    wire [71:0]d1_71__N_418;
    wire [71:0]d2_71__N_490;
    wire [71:0]d3_71__N_562;
    wire [71:0]d4_71__N_634;
    wire [71:0]d5_71__N_706;
    
    wire n15854, n168;
    wire [71:0]d6_71__N_1459;
    wire [71:0]d7_71__N_1531;
    wire [71:0]d8_71__N_1603;
    wire [71:0]d9_71__N_1675;
    
    wire n165, n183, n180_adj_2763, n177_adj_2764, n174_adj_2765, 
        n171_adj_2766, n168_adj_2767, n165_adj_2768, n162, n159, n156, 
        n153, n150, n147, n144, n141, n138, n135, n132, n129, 
        n126, n123, n120, n117, n114, n111, n108, n105, n102, 
        n99, n96, n93, n90_adj_2769, n87_adj_2770, n84_adj_2771, 
        n81_adj_2772, n78_adj_2773, n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, 
        n274, n271, n268, n265, n262, n259, n256, n253, n250, 
        n247, n244, n241, n238, n235, n232, n229, n226, n223, 
        n220, n217, n214, n211, n208, n205, n202, n199, n196, 
        n193, n190, n187, n184, n181, n178, n175, n172, n169, 
        n166, n163, n160, n157, n154, n151, n148, n145, n142, 
        n139, n136, n133, n130;
    wire [71:0]d_tmp_adj_5665;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(30[26:31])
    wire [71:0]d_d_tmp_adj_5666;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(30[33:40])
    wire [71:0]d1_adj_5667;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(35[26:28])
    wire [71:0]d2_adj_5668;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(36[26:28])
    wire [71:0]d3_adj_5669;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(37[26:28])
    wire [71:0]d4_adj_5670;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(38[26:28])
    wire [71:0]d5_adj_5671;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(39[26:28])
    wire [71:0]d6_adj_5672;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(43[26:28])
    wire [71:0]d_d6_adj_5673;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(43[30:34])
    wire [71:0]d7_adj_5674;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(44[26:28])
    wire [71:0]d_d7_adj_5675;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(44[30:34])
    wire [71:0]d8_adj_5676;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(45[26:28])
    wire [71:0]d_d8_adj_5677;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(45[30:34])
    wire [71:0]d9_adj_5678;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(46[26:28])
    wire [71:0]d_d9_adj_5679;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(46[30:34])
    wire [71:0]d10_adj_5680;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(47[26:29])
    
    wire n16053, n162_adj_3854, n159_adj_3855;
    wire [15:0]count_adj_5682;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(50[14:19])
    wire [71:0]d1_71__N_418_adj_5683;
    wire [71:0]d2_71__N_490_adj_5684;
    wire [71:0]d3_71__N_562_adj_5685;
    wire [71:0]d4_71__N_634_adj_5686;
    wire [71:0]d5_71__N_706_adj_5687;
    
    wire n16209, n16208, n16207, n16206, n16205, n16204, n16203, 
        n16202, n16201, n16200, n16199, n16198, n16197, n321, 
        n318, n315, n312, n309, n306, n303, n300, n297, n294, 
        n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255;
    wire [71:0]d6_71__N_1459_adj_5699;
    wire [71:0]d7_71__N_1531_adj_5700;
    wire [71:0]d8_71__N_1603_adj_5701;
    wire [71:0]d9_71__N_1675_adj_5702;
    
    wire n156_adj_4520, n15838, n15837, n15836, n15835, n15834, 
        n15833, n15832, n15831, n15830, n15829, n15827, n15826, 
        n15825, n15824, n15823, n15822, n15821, n15820, n15819, 
        n15818, n15817, n15816, n15815, n15814, n15813, n15812, 
        n15811, n15810;
    wire [71:0]d_out_11__N_1819_adj_5705;
    
    wire n252, n249, n246, n243, n240, n237, n234, n231, n228, 
        n225, n222, n219, n216, n213, n210, n207, n204, n201, 
        n198, n195, n192, n189, n186, n183_adj_4521, n180_adj_4522, 
        n177_adj_4523, n174_adj_4524, n171_adj_4525, n168_adj_4526, 
        n165_adj_4527, n162_adj_4528, n159_adj_4529, n156_adj_4530, 
        n153_adj_4531, n150_adj_4532, n147_adj_4533, n144_adj_4534, 
        n141_adj_4535, n138_adj_4536, n135_adj_4537, n132_adj_4538, 
        n183_adj_4539, n153_adj_4540, n150_adj_4541, n147_adj_4542, 
        n144_adj_4543, n141_adj_4544, n138_adj_4545, n135_adj_4546, 
        n132_adj_4547, n129_adj_4548, n126_adj_4549, n123_adj_4550, 
        n120_adj_4551, n117_adj_4552, n114_adj_4553, n111_adj_4554, 
        n108_adj_4555, n15912, n105_adj_4556, n102_adj_4557, n99_adj_4558, 
        n96_adj_4559, n93_adj_4560, n16052, n90_adj_4561, n87_adj_4562, 
        n84_adj_4563, n81_adj_4564, n78_adj_4565, n16051, n16050, 
        n16049, n16048, n16047, n16046, n16045, n16044, n11_adj_4566, 
        n15914, n16043, n16042, n16041, n16040;
    wire [9:0]counter;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(7[11:18])
    wire [11:0]DataInReg;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(10[12:21])
    
    wire n16039;
    wire [11:0]DataInReg_11__N_1856;
    
    wire n15806, n15805;
    wire [31:0]ISquare;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(24[14:21])
    
    wire n4_adj_4567, n3_adj_4568, n2_adj_4569;
    wire [23:0]MultResult1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(30[22:33])
    wire [23:0]MultResult2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(35[22:33])
    
    wire n22_adj_4570, n21_adj_4571, n20_adj_4572, n19_adj_4573, n18_adj_4574, 
        n17_adj_4575, n16_adj_4576, n16038, n2327, n16037, n15910, 
        n2326, n15_adj_4577, n16036, n2325, n2324, n14_adj_4578, 
        n209, n2323, n2322, n13_adj_4579, n2321, n2320, n37_adj_4580, 
        n36_adj_4581, n35_adj_4582, n34_adj_4583, n33_adj_4584, n32_adj_4585, 
        n31_adj_4586, n30_adj_4587, n29_adj_4588, n28_adj_4589, n27_adj_4590, 
        n26_adj_4591, n12_adj_4592, n25_adj_4593, n2319, n24_adj_4594, 
        n23_adj_4595, n22_adj_4596, n21_adj_4597, n20_adj_4598, n19_adj_4599, 
        n18_adj_4600, n17_adj_4601, n16_adj_4602, n15_adj_4603, n14_adj_4604, 
        n13_adj_4605, n12_adj_4606, n11_adj_4607, n10_adj_4608, n9_adj_4609, 
        n8_adj_4610, n7_adj_4611, n6_adj_4612, n5_adj_4613, n4_adj_4614, 
        n3_adj_4615, n2_adj_4616;
    wire [17:0]d_out_d_11__N_1874;
    
    wire d_out_d_11__N_1873, n11_adj_4617, n2317, n2316, n37_adj_4618, 
        n36_adj_4619, n35_adj_4620, n34_adj_4621, n33_adj_4622, n32_adj_4623, 
        n31_adj_4624;
    wire [17:0]d_out_d_11__N_1876;
    
    wire d_out_d_11__N_1875, n10_adj_4625, n30_adj_4626, n2315, n29_adj_4627, 
        n28_adj_4628, n27_adj_4629, n26_adj_4630, n25_adj_4631, n24_adj_4632, 
        n23_adj_4633, n22_adj_4634, n21_adj_4635, n20_adj_4636, n19_adj_4637, 
        n18_adj_4638, n17_adj_4639, n16_adj_4640, n15_adj_4641, n14_adj_4642, 
        n13_adj_4643, n2314, n12_adj_4644, n11_adj_4645, n10_adj_4646, 
        n9_adj_4647, n8_adj_4648, n7_adj_4649, n6_adj_4650, n5_adj_4651, 
        n4_adj_4652, n3_adj_4653, n2_adj_4654;
    wire [17:0]d_out_d_11__N_1878;
    
    wire d_out_d_11__N_1877, n9_adj_4655, n2313, n2312, n37_adj_4656, 
        n36_adj_4657;
    wire [17:0]d_out_d_11__N_1880;
    
    wire d_out_d_11__N_1879, n8_adj_4658, n35_adj_4659, n2311, n34_adj_4660, 
        n33_adj_4661, n32_adj_4662, n31_adj_4663, n30_adj_4664, n29_adj_4665, 
        n28_adj_4666, n27_adj_4667, n26_adj_4668, n25_adj_4669, n24_adj_4670, 
        n23_adj_4671, n22_adj_4672, n21_adj_4673, n20_adj_4674, n19_adj_4675, 
        n18_adj_4676, n2310, n17_adj_4677, n16_adj_4678, n15_adj_4679, 
        n14_adj_4680, n13_adj_4681, n9_adj_4682, n10_adj_4683, n11_adj_4684, 
        n12_adj_4685, n8_adj_4686;
    wire [17:0]d_out_d_11__N_1882;
    
    wire n7_adj_4687, n37_adj_4688, n6_adj_4689, n5_adj_4690, n4_adj_4691, 
        n3_adj_4692, n2_adj_4693, n36_adj_4694, n35_adj_4695, n34_adj_4696, 
        n33_adj_4697;
    wire [17:0]d_out_d_11__N_1884;
    
    wire n15877, n15853, n15852, n15851, n15850, n3691, n15859, 
        n15860, n15879, n15862, n15864, n15865, n15866, n15872, 
        n15873, n15874, n3677, n3676;
    wire [17:0]d_out_d_11__N_1886;
    
    wire n15878, n15858, n15880, n15884, n15881, n15882, n15883, 
        n15875, n15885, n15886, n15887, n15888, n15896, n15876, 
        n3659, n3656, n15894, n15892, n15895, n14928, n15846, 
        n15845, n15844;
    wire [17:0]d_out_d_11__N_1888;
    
    wire n15843, n37_adj_4698, n36_adj_4699;
    wire [17:0]d_out_d_11__N_1890;
    
    wire n35_adj_4700, n34_adj_4701, n33_adj_4702, n32_adj_4703, n31_adj_4704, 
        n30_adj_4705, n29_adj_4706, n28_adj_4707, n27_adj_4708, n26_adj_4709, 
        n25_adj_4710, n24_adj_4711, n23_adj_4712, n22_adj_4713, n21_adj_4714, 
        n20_adj_4715, n19_adj_4716, n18_adj_4717, n17_adj_4718, n16_adj_4719, 
        n15_adj_4720, n14_adj_4721, n13_adj_4722, n12_adj_4723, n11_adj_4724, 
        n10_adj_4725, n9_adj_4726, n8_adj_4727, n7_adj_4728, n6_adj_4729, 
        n15909;
    wire [17:0]d_out_d_11__N_1892;
    
    wire n912, n913, n914, n915, n916, n917, n918, n919, n920, 
        n921, n922, n923, n924, n925, n926, n927, n5_adj_4730;
    wire [17:0]d_out_d_11__N_2353;
    
    wire n16196, n16035, n16195, n16034, n16194;
    wire [17:0]d_out_d_11__N_2335;
    
    wire n16033, n2330, n16032, n16031, n16030, n16029, n2332, 
        n16028, n16027, n16026, n2336, n15804, n16_adj_4731, n16193, 
        n16192, n16188, n16187, n16186, n16185, n16184, n15803, 
        n15802, n2334, n2335, n16183, n16182, n16181, n16180, 
        n16179, n16178, n16177, n16176, n16175, n16174, n16173, 
        n15908, n15801, n15907, n16025, n16024, n16023, n16022, 
        n16021, n2333, n16172, n16171, n16170, n16169, n16168, 
        n16167, n16166, n16165, n16164, n15800, n15799, n15798, 
        n16019, n16018, n16017, n16016, n16163, n16162, n16161, 
        n16160, n16159, n15797, n15796, n15795, n15792, n15791, 
        n15790, n15789, n15788, n15787, n15786, n15785, n15784, 
        n15783, n15782, n15781, n15780, n15779, n15778, n16015, 
        n16014, n17628, n16013, n16012, n10_adj_4732, n183_adj_4733, 
        n16011, n180_adj_4734, n177_adj_4735, n174_adj_4736, n16158, 
        n15842, n2369, n2368, n2367, n2366, n2365, n2363, n2362, 
        n2361, n2360, n2359, n2358, n2356, n2355, n2354, n2352, 
        n2350, n2349, n2559, n2558, n16157, n2555, n16156, n16155, 
        n2549, n2548, n15841, n2541, n15840, n2530, n16154, n16153, 
        n16152, n2520, n16151, clk_80mhz_enable_1470, n16150, n2514, 
        n2513, n171_adj_4737, n168_adj_4738, n16010, n16009, n16008, 
        n16007, n16006, n16005, n16004, n16003, n16002, n15998, 
        n15997, n15996, n15995, n15906, n2636, n16149, n15994, 
        n15993, n16148, n165_adj_4739, n15777, n162_adj_4740, n159_adj_4741, 
        n156_adj_4742, n17625, n17751, n63, n64, n17642, n66, 
        n67, n153_adj_4743, n150_adj_4744, n17750, n147_adj_4745, 
        n144_adj_4746, n15992, n16147, n141_adj_4747, n138_adj_4748, 
        n16146, n16145, n16144, n135_adj_4749, n2348, n2347, n2346, 
        n2345, n2344, n2343, n2342, n2341, n2340, n2339, n2338, 
        n2337, n132_adj_4750, n16143, n16142, n16141, n15_adj_4751, 
        n14_adj_4752, n13_adj_4753, n12_adj_4754, n11_adj_4755, n10_adj_4756, 
        n9_adj_4757, n8_adj_4758, n7_adj_4759, n6_adj_4760, n5_adj_4761, 
        n4_adj_4762, n3_adj_4763, n2_adj_4764, n15991, n129_adj_4765, 
        n126_adj_4766, n123_adj_4767, n16140, n16139, n16138, n16137, 
        n16136, n16135, n16134, n16133, n2571, clk_80mhz_enable_1408, 
        n16132, n37_adj_4768, n16131, n36_adj_4769, n35_adj_4770, 
        n34_adj_4771, n33_adj_4772, n32_adj_4773, n16130, n31_adj_4774, 
        n30_adj_4775, n29_adj_4776, n28_adj_4777, n27_adj_4778, n26_adj_4779, 
        n25_adj_4780, n24_adj_4781, n15990, n15989, n16129, n120_adj_4782, 
        n117_adj_4783, n114_adj_4784, n111_adj_4785, n2823, n16128, 
        n2328, n108_adj_4786, n105_adj_4787, n16084, n102_adj_4788, 
        n99_adj_4789, n15988, n96_adj_4790, n15776, n17_adj_4791, 
        n15905, n18_adj_4792, n35_adj_4793, n34_adj_4794, n33_adj_4795, 
        n32_adj_4796, n31_adj_4797, n30_adj_4798, n29_adj_4799, n28_adj_4800, 
        n27_adj_4801, n26_adj_4802, n25_adj_4803, n24_adj_4804, n23_adj_4805, 
        n22_adj_4806, n21_adj_4807, n20_adj_4808, n19_adj_4809, n36_adj_4810, 
        n37_adj_4811, n24_adj_4812, n15987, n15986, n93_adj_4813, 
        n23_adj_4814, n22_adj_4815, n21_adj_4816, n20_adj_4817, n19_adj_4818, 
        n18_adj_4819, n17_adj_4820, n16_adj_4821, n15_adj_4822, n14_adj_4823, 
        n13_adj_4824, n12_adj_4825, n11_adj_4826, n10_adj_4827, n9_adj_4828, 
        n8_adj_4829, n7_adj_4830, n6_adj_4831, n5_adj_4832, n4_adj_4833, 
        n3_adj_4834, n2_adj_4835, n23_adj_4836, n16127, cout_adj_4837, 
        n78_adj_4838, n81_adj_4839, n84_adj_4840, n87_adj_4841, n90_adj_4842, 
        n93_adj_4843, n96_adj_4844, n99_adj_4845, n102_adj_4846, n105_adj_4847, 
        n108_adj_4848, n111_adj_4849, n114_adj_4850, n117_adj_4851, 
        n120_adj_4852, n123_adj_4853, n126_adj_4854, n129_adj_4855, 
        n132_adj_4856, n135_adj_4857, n138_adj_4858, n141_adj_4859, 
        n144_adj_4860, n147_adj_4861, n150_adj_4862, n153_adj_4863, 
        n156_adj_4864, n159_adj_4865, n162_adj_4866, n165_adj_4867, 
        n168_adj_4868, n171_adj_4869, n174_adj_4870, n177_adj_4871, 
        n180_adj_4872, n183_adj_4873, n78_adj_4874, n81_adj_4875, n84_adj_4876, 
        n87_adj_4877, n90_adj_4878, n93_adj_4879, n96_adj_4880, n99_adj_4881, 
        n102_adj_4882, n105_adj_4883, n108_adj_4884, n111_adj_4885, 
        n114_adj_4886, n117_adj_4887, n120_adj_4888, n78_adj_4889, n81_adj_4890, 
        n84_adj_4891, n87_adj_4892, n90_adj_4893, n93_adj_4894, n96_adj_4895, 
        n99_adj_4896, n102_adj_4897, n105_adj_4898, n108_adj_4899, n111_adj_4900, 
        n114_adj_4901, n117_adj_4902, n120_adj_4903, n123_adj_4904, 
        n126_adj_4905, n129_adj_4906, n132_adj_4907, n135_adj_4908, 
        n138_adj_4909, n141_adj_4910, n144_adj_4911, n147_adj_4912, 
        n150_adj_4913, n153_adj_4914, n156_adj_4915, n159_adj_4916, 
        n162_adj_4917, n165_adj_4918, n168_adj_4919, n171_adj_4920, 
        n174_adj_4921, n177_adj_4922, n180_adj_4923, n183_adj_4924, 
        n78_adj_4925, n81_adj_4926, n84_adj_4927, n87_adj_4928, n90_adj_4929, 
        n93_adj_4930, n96_adj_4931, n99_adj_4932, n102_adj_4933, n105_adj_4934, 
        n108_adj_4935, n111_adj_4936, n114_adj_4937, n117_adj_4938, 
        n120_adj_4939, n123_adj_4940, n126_adj_4941, n129_adj_4942, 
        n132_adj_4943, n135_adj_4944, n138_adj_4945, n141_adj_4946, 
        n144_adj_4947, n147_adj_4948, n150_adj_4949, n153_adj_4950, 
        n156_adj_4951, n159_adj_4952, n162_adj_4953, n165_adj_4954, 
        n168_adj_4955, n171_adj_4956, n174_adj_4957, n177_adj_4958, 
        n180_adj_4959, n183_adj_4960, n78_adj_4961, n81_adj_4962, n84_adj_4963, 
        n87_adj_4964, n90_adj_4965, n93_adj_4966, n96_adj_4967, n99_adj_4968, 
        n102_adj_4969, n105_adj_4970, n108_adj_4971, n111_adj_4972, 
        n114_adj_4973, n117_adj_4974, n120_adj_4975, n123_adj_4976, 
        n126_adj_4977, n129_adj_4978, n132_adj_4979, n135_adj_4980, 
        n138_adj_4981, n141_adj_4982, n144_adj_4983, n147_adj_4984, 
        n150_adj_4985, n153_adj_4986, n156_adj_4987, n159_adj_4988, 
        n162_adj_4989, n165_adj_4990, n168_adj_4991, n171_adj_4992, 
        n174_adj_4993, n177_adj_4994, n180_adj_4995, n183_adj_4996, 
        n134, n137, n140, n143, n146, n149, n152, n155, n158, 
        n161, n164, n167, n170, n173, n176, n179, n182, n185, 
        n188, n191, n194, n197, n200, n203, n206, n209_adj_4997, 
        n212, n215, n218, n221, n224, n227, n230, n233, n236, 
        n239, n242, n245, n248, n251, n254, n257, n260, n263, 
        n266, n269, n272, n275, n278, n281, n284, n287, n290, 
        n293, n296, n299, n302, n305, n308, n311, n314, n317, 
        n320, n323, n15775, n15771, n15770, n15769, n15768, n15767, 
        n15766, n15765, cout_adj_4998, cout_adj_4999, cout_adj_5000, 
        n78_adj_5001, n81_adj_5002, n84_adj_5003, n87_adj_5004, n90_adj_5005, 
        n93_adj_5006, n96_adj_5007, n99_adj_5008, n102_adj_5009, n105_adj_5010, 
        n108_adj_5011, n111_adj_5012, n114_adj_5013, n117_adj_5014, 
        n120_adj_5015, n123_adj_5016, n126_adj_5017, n129_adj_5018, 
        n132_adj_5019, n135_adj_5020, n138_adj_5021, n141_adj_5022, 
        n144_adj_5023, n147_adj_5024, n150_adj_5025, n153_adj_5026, 
        n156_adj_5027, n159_adj_5028, n162_adj_5029, n165_adj_5030, 
        n168_adj_5031, n171_adj_5032, n174_adj_5033, n177_adj_5034, 
        n180_adj_5035, n183_adj_5036, n78_adj_5037, n81_adj_5038, n84_adj_5039, 
        n87_adj_5040, n90_adj_5041, n93_adj_5042, n96_adj_5043, n99_adj_5044, 
        n102_adj_5045, n105_adj_5046, n108_adj_5047, n111_adj_5048, 
        n114_adj_5049, n117_adj_5050, n120_adj_5051, n78_adj_5052, n81_adj_5053, 
        n84_adj_5054, n87_adj_5055, n90_adj_5056, n93_adj_5057, n96_adj_5058, 
        n99_adj_5059, n102_adj_5060, n105_adj_5061, n108_adj_5062, n111_adj_5063, 
        n114_adj_5064, n117_adj_5065, n120_adj_5066, n123_adj_5067, 
        n126_adj_5068, n129_adj_5069, n132_adj_5070, n135_adj_5071, 
        n138_adj_5072, n141_adj_5073, n144_adj_5074, n147_adj_5075, 
        n150_adj_5076, n153_adj_5077, n156_adj_5078, n159_adj_5079, 
        n162_adj_5080, n165_adj_5081, n168_adj_5082, n171_adj_5083, 
        n174_adj_5084, n177_adj_5085, n180_adj_5086, n183_adj_5087, 
        cout_adj_5088, n15764, n15763, n15762, n15761, n15760, n15759, 
        n15758, n15757, n15756, n15755, n15754, n15753, n15752, 
        n15751, n15750, n15749, n15748, n15747, n15746, n15745, 
        n15744, n15743, n15742, n15741, n15740, n15739, n15738, 
        n15737, n15736, n15735, n15734, n15733, n15732, n15731, 
        n15730, n15729, cout_adj_5089, n78_adj_5090, n81_adj_5091, 
        n84_adj_5092, n87_adj_5093, n90_adj_5094, n93_adj_5095, n96_adj_5096, 
        n99_adj_5097, n102_adj_5098, n105_adj_5099, n108_adj_5100, n111_adj_5101, 
        n114_adj_5102, n117_adj_5103, n120_adj_5104, n123_adj_5105, 
        n126_adj_5106, n129_adj_5107, n132_adj_5108, n135_adj_5109, 
        n138_adj_5110, n141_adj_5111, n144_adj_5112, n147_adj_5113, 
        n150_adj_5114, n153_adj_5115, n156_adj_5116, n159_adj_5117, 
        n162_adj_5118, n165_adj_5119, n168_adj_5120, n171_adj_5121, 
        n174_adj_5122, n177_adj_5123, n180_adj_5124, n183_adj_5125, 
        cout_adj_5126, cout_adj_5127, cout_adj_5128, n36_adj_5129, n39, 
        n42, n45, n48, n51, n54, n57, n60, n63_adj_5130, n66_adj_5131, 
        n69, n72, n75, n78_adj_5132, n81_adj_5133, cout_adj_5134, 
        cout_adj_5135, cout_adj_5136, cout_adj_5137, n36_adj_5138, n39_adj_5139, 
        n42_adj_5140, n45_adj_5141, n48_adj_5142, n51_adj_5143, n54_adj_5144, 
        n57_adj_5145, n60_adj_5146, n63_adj_5147, n66_adj_5148, n69_adj_5149, 
        n72_adj_5150, n75_adj_5151, n78_adj_5152, n81_adj_5153, n76, 
        n79, n82, n85, n88, n91, n94, n97, n100, n103, n106, 
        n109, n112, n115, n118, n54_adj_5154, n57_adj_5155, n60_adj_5156, 
        n63_adj_5157, n66_adj_5158, n69_adj_5159, n72_adj_5160, n75_adj_5161, 
        n78_adj_5162, n81_adj_5163, n84_adj_5164, n87_adj_5165, n90_adj_5166, 
        n93_adj_5167, n96_adj_5168, n99_adj_5169, n102_adj_5170, n105_adj_5171, 
        n108_adj_5172, n111_adj_5173, n114_adj_5174, n117_adj_5175, 
        n120_adj_5176, n123_adj_5177, n126_adj_5178, cout_adj_5179, 
        n78_adj_5180, n81_adj_5181, n84_adj_5182, n87_adj_5183, n90_adj_5184, 
        n93_adj_5185, n96_adj_5186, n99_adj_5187, n102_adj_5188, n105_adj_5189, 
        n108_adj_5190, n111_adj_5191, n114_adj_5192, n117_adj_5193, 
        n120_adj_5194, n123_adj_5195, n126_adj_5196, n129_adj_5197, 
        n132_adj_5198, n135_adj_5199, n138_adj_5200, n141_adj_5201, 
        n144_adj_5202, n147_adj_5203, n150_adj_5204, n153_adj_5205, 
        n156_adj_5206, n159_adj_5207, n162_adj_5208, n165_adj_5209, 
        n168_adj_5210, n171_adj_5211, n174_adj_5212, n177_adj_5213, 
        n180_adj_5214, n183_adj_5215, cout_adj_5216, cout_adj_5217, 
        n78_adj_5218, n81_adj_5219, n84_adj_5220, n87_adj_5221, n90_adj_5222, 
        n93_adj_5223, n96_adj_5224, n99_adj_5225, n102_adj_5226, n105_adj_5227, 
        n108_adj_5228, n111_adj_5229, n114_adj_5230, n117_adj_5231, 
        n120_adj_5232, n123_adj_5233, n126_adj_5234, n129_adj_5235, 
        n132_adj_5236, n135_adj_5237, n138_adj_5238, n141_adj_5239, 
        n144_adj_5240, n147_adj_5241, n150_adj_5242, n153_adj_5243, 
        n156_adj_5244, n159_adj_5245, n162_adj_5246, n165_adj_5247, 
        n168_adj_5248, n171_adj_5249, n174_adj_5250, n177_adj_5251, 
        n180_adj_5252, n183_adj_5253, cout_adj_5254, n16126, n16083, 
        n12132, n16125, n16082, n12134, n16124, n12136, n16123, 
        n12108, n12138, n16122, n16081, n12140, n16121, n16080, 
        n12142, n16120, n16079, n12144, n16119, n16078, n12146, 
        n16118, n16077, n16059, n16075, n16074, n16073, n51_adj_5255, 
        n54_adj_5256, n57_adj_5257, n60_adj_5258, n63_adj_5259, n15985, 
        n66_adj_5260, n69_adj_5261, n15984, n72_adj_5262, n75_adj_5263, 
        n15911, n78_adj_5264, n81_adj_5265, n16072, n84_adj_5266, 
        n87_adj_5267, n16071, n90_adj_5268, n15983, n15982, n16067, 
        n15981, n15978, n15977, n16066, n15976, n15975, n12148, 
        n12023, n12021, n12019, n12013, n12011, n17638, n12007, 
        n12003, n12001, n11999, n11997, n11995, n11993, n11989, 
        n11987, n11985, n11983, n11981, n11979, n78_adj_5269, n11977, 
        n81_adj_5270, n11975, n84_adj_5271, n11973, n87_adj_5272, 
        n11971, n90_adj_5273, n93_adj_5274, n96_adj_5275, n11967, 
        n99_adj_5276, n11965, n102_adj_5277, n11963, n105_adj_5278, 
        n11961, n108_adj_5279, n11959, n111_adj_5280, n11957, n114_adj_5281, 
        n117_adj_5282, n120_adj_5283, n11953, n123_adj_5284, n126_adj_5285, 
        n129_adj_5286, n11949, n132_adj_5287, n135_adj_5288, n138_adj_5289, 
        n11945, n141_adj_5290, n11943, n144_adj_5291, n147_adj_5292, 
        n150_adj_5293, n153_adj_5294, n16399, n156_adj_5295, n11937, 
        n159_adj_5296, n11935, n162_adj_5297, n11933, n165_adj_5298, 
        n168_adj_5299, n16398, n171_adj_5300, n11929, n174_adj_5301, 
        n11927, n177_adj_5302, n12511, n180_adj_5303, n183_adj_5304, 
        n16397, n16396, n16395, n16394, n16393, n16812, n16117, 
        n12378, n78_adj_5305, n81_adj_5306, n84_adj_5307, n87_adj_5308, 
        n90_adj_5309, n93_adj_5310, n96_adj_5311, n99_adj_5312, n102_adj_5313, 
        n105_adj_5314, n108_adj_5315, n111_adj_5316, n114_adj_5317, 
        n117_adj_5318, n120_adj_5319, n123_adj_5320, n126_adj_5321, 
        n129_adj_5322, n132_adj_5323, n135_adj_5324, n15974, n138_adj_5325, 
        n15973, n141_adj_5326, n15972, n144_adj_5327, n15971, n147_adj_5328, 
        n15970, n150_adj_5329, n15969, n153_adj_5330, n15968, n156_adj_5331, 
        n15967, n159_adj_5332, n15966, n162_adj_5333, n15965, n165_adj_5334, 
        n15964, n168_adj_5335, n15963, n171_adj_5336, n15962, n174_adj_5337, 
        n15961, n177_adj_5338, n180_adj_5339, n16115, n183_adj_5340, 
        n16387, n15867, n16060, n16386, n16385, n16384, n15957, 
        n16114, n16113, n16383, n15956, n16382, n16112, n16111, 
        n15955, n16381, n16110, n15857, n16109, n16380, n16108, 
        n15954, n16379, n16107, n15953, n16106, n11690, n16105, 
        n15952, n16104, n15863, n16103, n15951, n16373, clk_80mhz_enable_1471, 
        n16102, n16101, n15950, n16372, n15949, n16371, n16370, 
        n16100, n15889, n16369, n15948, n16099, n15947, n16098, 
        n16368, n16367, n15891, n16094, n15946, n16366, n15728, 
        n15727, n15726, n15725, n15724, n15723, n15722, n15721, 
        n15720, n15719, n15718, n15717, n15716, n15715, n15714, 
        n15713, cout_adj_5341, n16093, n15712, n16065, n15945, n16364, 
        n16363, n15904, n16362, n16092, n16361, n16091, n15944, 
        n15861, n16360, n16064, n16090, n15903, n16359, n15943, 
        n16358, n15942, n16357, n16089, n16088, n15902, n16356, 
        n16355, n15941, n15711, n15940, n15938, n15937, n15936, 
        n15935, n15934, n15933, n15932, n15931, n15930, n15929, 
        n15928, n15927, n15926, n16354, n16353, n15925, n16087, 
        n16352, n16351, n16350, n16086, n15924, n15897, n15923, 
        n15922, n15921, n15919, n15918, n15917, n15916, n15915, 
        n16349, n16348, n16347, n16346, n16345, n16344, n16343, 
        n16070, n16342, n16063, n16341, n17304, n78_adj_5342, n81_adj_5343, 
        n84_adj_5344, n87_adj_5345, n90_adj_5346, n93_adj_5347, n96_adj_5348, 
        n99_adj_5349, n102_adj_5350, n16340, n105_adj_5351, n108_adj_5352, 
        n16339, n111_adj_5353, n114_adj_5354, n117_adj_5355, n120_adj_5356, 
        n16338, n123_adj_5357, n126_adj_5358, n16337, n129_adj_5359, 
        n132_adj_5360, n135_adj_5361, n16336, n138_adj_5362, n15893, 
        n141_adj_5363, n16335, n144_adj_5364, n147_adj_5365, n16334, 
        n150_adj_5366, n153_adj_5367, n16333, n156_adj_5368, n16062, 
        n159_adj_5369, n162_adj_5370, n165_adj_5371, n168_adj_5372, 
        n15898, n171_adj_5373, n174_adj_5374, n177_adj_5375, n180_adj_5376, 
        n16328, n183_adj_5377, n16327, n16326, n16325, n16061, n16324, 
        n16323, n16322, n16321, n16315, n16314, n16313, n16312, 
        n16311, n16310, n16069, n16309, n16308, n16307, n16068, 
        n16301, n16300, n16299, n16298, n17637, n16297, n16296, 
        n15856, n16290, n15855, n16289, n16288, n16287, n16286, 
        n16285, n16284, n16283, n16282, n16085, n15710, n15709, 
        n15708, n15707, n15706, n15705, n15704, n15703, n15702, 
        n15701, n15700, n15699, n15698, n15697, n15696, n15695, 
        n15694, n15693, n15692, n15691, n15690, n15689, n15688, 
        n15687, n15686, n15685, n15684, n15683, n15682, n15681, 
        n15680, n15679, n15678, n15677, n15676, n15675, n15674, 
        n15673, n15672, n15671, n15670, n15669, n15668, n15667, 
        n15666, n15665, n15664, n15663, n15662, n15661, n15660, 
        n15659, n15658, n15657, n15656, n15655, n15653, n15652, 
        n15651, n15650, n15649, n15648, n15647, n15646, n15645, 
        n15644, n15643, n15642, n15641, n15640, n15639, n15638, 
        n15637, n15636, n15635, n15634, n15633, n15632, n15631, 
        n15630, n15629, n15628, n15627, n15626, n52, n15625, n55, 
        n15624, n58, n15623, n61, n15621, n64_adj_5378, n15620, 
        n67_adj_5379, n15619, n70, n15618, n73, n15617, n76_adj_5380, 
        n15616, n79_adj_5381, n15615, n82_adj_5382, n15614, n85_adj_5383, 
        n15613, n15612, n15611, n15610, n15609, n15608, n15607, 
        n15606, n15605, n15604, n15603, n15602, n15601, n15600, 
        n15599, n15598, n15597, n15596, n15595, n15594, n15593, 
        n15591, n15590, n15589, n15588, n15587, n15586, n15585, 
        n15584, n15583, n15582, n15581, n15580, n15579, n15578, 
        n15577, n15576, n15575, n15574, n15570, n15569, n15568, 
        n15567, n15566, n15565, n15564, n15563, n15562, n15561, 
        n15560, n15559, n15558, n15557, n15556, n15555, n15554, 
        n15553, n15551, n15550, n15549, n15548, n15547, n15546, 
        n15545, n15544, n15543, n15542, n15541, n15540, n15539, 
        n15538, n15537, n15536, n15535, n15534, n15530, n15529, 
        n15528, n15527, n15526, n15525, n15523, n15522, n15521, 
        n15520, n15519, n15518, n15517, n15516, n15515, n15514, 
        n15513, n15512, n15511, n15510, n15509, n15508, n15507, 
        n15506, n15505, n15504, n15503, n15502, n15501, n15500, 
        n15499, n15498, n15497, n15496, n15495, n15494, n15493, 
        n15492, n15491, n15490, n15489, n15488, n15487, n15486, 
        n15485, n15484, n15483, n15482, n15481, n15480, n15479, 
        n15478, n15477, n15476, n15475, n15473, n15472, n15471, 
        n15470, n15469, n15468, n15467, n15466, n15465, n15464, 
        n15463, n15462, n15461, n15460, n15459, n15458, n15457, 
        n15456, n15452, n15451, n15450, n15449, n15448, n15447, 
        n15446, n15445, n15444, n15443, n15442, n15441, n78_adj_5384, 
        n15440, n81_adj_5385, n15439, n84_adj_5386, n15438, n87_adj_5387, 
        n15437, n90_adj_5388, n15436, n93_adj_5389, n15435, n96_adj_5390, 
        n99_adj_5391, n15433, n102_adj_5392, n15432, n105_adj_5393, 
        n15431, n108_adj_5394, n15430, n111_adj_5395, n15429, n114_adj_5396, 
        n15428, n117_adj_5397, n15427, n120_adj_5398, n15426, n123_adj_5399, 
        n15425, n126_adj_5400, n15424, n129_adj_5401, n15423, n132_adj_5402, 
        n15422, n135_adj_5403, n15421, n138_adj_5404, n15420, n141_adj_5405, 
        n15419, n144_adj_5406, n15418, n147_adj_5407, n15417, n150_adj_5408, 
        n15416, n153_adj_5409, n156_adj_5410, n159_adj_5411, n15412, 
        n162_adj_5412, n15411, n165_adj_5413, n15410, n168_adj_5414, 
        n15409, n171_adj_5415, n15408, n174_adj_5416, n15407, n177_adj_5417, 
        n15406, n180_adj_5418, n15405, n183_adj_5419, n15404, n15403, 
        n15402, n15401, n15400, n15399, n15398, n15397, n15396, 
        n15395, n15394, n15393, n15392, n15391, n15390, n15389, 
        n15388, n15387, n15386, n15385, n15384, n15383, n15382, 
        n15381, n15380, n15379, n15378, n15377, n15375, n15374, 
        n15373, n15372, n15371, n15370, n15369, n15368, n15367, 
        n15366, n15365, n15364, n15363, n15362, n15361, n15360, 
        n15359, n15358, n15353, n15352, n15351, n15350, n15349, 
        n15348, n15347, n15346, n15345, n15344, n15343, n15342, 
        n15341, n15340, n15339, n15338, n15337, n15336, n15331, 
        n15330, n15329, n15328, n15327, n15326, n15325, n15324, 
        n15323, n15322, n15321, n15320, n15319, n15318, n15317, 
        n15316, n15315, n15314, n15309, n15308, n15307, n15306, 
        n15305, n15304, n15303, n15302, n15301, n15300, n15299, 
        n15298, n15297, n15296, n15295, n15294, n15293, n15292, 
        n15288, n15287, cout_adj_5420, n15286, n15285, n15284, n15283, 
        n15282, n15281, n15280, n15279, n15278, n15277, n15276, 
        n15275, n15274, n15273, n15272, n15271, n15270, n15269, 
        n15268, n15267, n15266, n15265, n15264, n15263, n15262, 
        n15261, n15260, n15259, n15258, n15257, n15256, n15255, 
        n15254, n15253, n15252, n15251, n15250, n15249, n15248, 
        n15247, n15246, n15245, n15244, n44, n47, n15243, n50, 
        n15242, n53, n15241, n56, n15240, n59, n15239, n62, 
        n15238, n65, n15237, n15236, n15235, n15234, n15233, n15232, 
        n15231, n15230, n15229, n15228, n15227, n15226, n15225, 
        n15224, n15223, n15222, n15221, n15220, n15219, n15218, 
        n15217, n15216, n15215, n15214, n15213, n15212, n15211, 
        n15210, n15209, n15208, n45_adj_5421, n15207, n48_adj_5422, 
        n15206, n51_adj_5423, n15205, n54_adj_5424, n15204, n57_adj_5425, 
        n15203, n60_adj_5426, n15202, n63_adj_5427, n15201, n66_adj_5428, 
        n15200, n69_adj_5429, n15199, n72_adj_5430, n15197, n75_adj_5431, 
        n15196, n78_adj_5432, n15195, n81_adj_5433, n15194, n84_adj_5434, 
        n15193, n87_adj_5435, n15192, n90_adj_5436, n15191, n15190, 
        n15189, n15188, n15187, n15186, n15185, n15184, n15183, 
        n15182, n15181, n15180, n15178, n15177, n15176, n15175, 
        n15174, n15173, n15172, n15171, n15170, n15169, n15168, 
        n15167, n15166, n15165, n15164, n15163, n15162, n15161, 
        n15159, n15158, n15157, n15156, n15155, n15154, n15153, 
        n15152, n15151, n15150, n15149, n15148, n15147, n15146, 
        n15145, n15144, n15143, n15142, n15140, n15139, n15138, 
        n15137, n15136, n15135, n15134, n15133, n15132, n15131, 
        n15130, n15129, n15128, n15127, n15126, n78_adj_5437, n15125, 
        n81_adj_5438, n84_adj_5439, n87_adj_5440, n90_adj_5441, n93_adj_5442, 
        n96_adj_5443, n99_adj_5444, n102_adj_5445, n105_adj_5446, n108_adj_5447, 
        n111_adj_5448, n114_adj_5449, n117_adj_5450, n120_adj_5451, 
        n123_adj_5452, n126_adj_5453, n129_adj_5454, n132_adj_5455, 
        n135_adj_5456, n138_adj_5457, n141_adj_5458, n144_adj_5459, 
        n147_adj_5460, n150_adj_5461, n153_adj_5462, n156_adj_5463, 
        n159_adj_5464, n162_adj_5465, n165_adj_5466, n168_adj_5467, 
        n171_adj_5468, n174_adj_5469, n177_adj_5470, n180_adj_5471, 
        n183_adj_5472, n15124, n15123, n15121, n15120, n15119, n15118, 
        n15117, n15116, n15115, n15114, n15113, n15112, n15111, 
        n15110, n15109, n15108, n15107, n15106, n15105, n15104, 
        n15102, n15101, n15100, n15099, n15098, n15097, n15096, 
        n15095, n15094, n15093, n15092, n15091, n15090, n15089, 
        n15088, n15087, n15086, n15085, n15084, n15083, n15082, 
        n15081, n15080, n15079, n15078, n15077, n15076, n15075, 
        n15074, n15073, n45_adj_5473, n15072, n48_adj_5474, n15071, 
        n51_adj_5475, n15070, n54_adj_5476, n15069, n57_adj_5477, 
        n15068, n60_adj_5478, n15067, n63_adj_5479, n15066, n66_adj_5480, 
        n15065, n69_adj_5481, n15064, n72_adj_5482, n15063, n75_adj_5483, 
        n15062, n78_adj_5484, n15061, n81_adj_5485, n15060, n84_adj_5486, 
        n15059, n87_adj_5487, n15058, n90_adj_5488, n15057, n15056, 
        n15055, n15054, n15053, n15052, n15051, n15050, n15049, 
        n15048, n15047, n15046, n15045, n15044, n15043, n15042, 
        n15041, n15040, n15039, n15038, n15037, n15036, n15035, 
        n15034, n15033, n15032, n15031, n15030, n15029, n15028, 
        n15027, n15026, n15025, n15024, n15023, n15022, n45_adj_5489, 
        n48_adj_5490, n15021, n51_adj_5491, n15020, n54_adj_5492, 
        n15019, n57_adj_5493, n15018, n60_adj_5494, n15017, n63_adj_5495, 
        n15016, n66_adj_5496, n15015, n69_adj_5497, n15014, n72_adj_5498, 
        n15013, n75_adj_5499, n15012, n78_adj_5500, n15011, n81_adj_5501, 
        n15010, n84_adj_5502, n15009, n87_adj_5503, n15008, n90_adj_5504, 
        n15007, n15006, n15005, n15004, n15003, n15002, n15001, 
        n15000, n14999, n14998, n14997, n14996, n14995, n14994, 
        n14993, n14992, n14991, n14990, n14989, n14988, n14987, 
        n14986, n14985, n14984, n14983, n14982, n14981, n14980, 
        n14979, n14978, n14977, n14976, n14975, n14974, n14973, 
        n14972, n14971, n14970, n14969, n14968, n45_adj_5505, n14967, 
        n48_adj_5506, n14966, n51_adj_5507, n14965, n54_adj_5508, 
        n14964, n57_adj_5509, n14963, n60_adj_5510, n14962, n63_adj_5511, 
        n14961, n66_adj_5512, n14960, n69_adj_5513, n14959, n72_adj_5514, 
        n14958, n75_adj_5515, n14957, n78_adj_5516, n81_adj_5517, 
        n14955, n84_adj_5518, n14954, n87_adj_5519, n14953, n90_adj_5520, 
        n14952, n14951, n14950, n14949, n14948, n14947, n14946, 
        n14945, n14944, n14943, n14942, n14941, n14940, n14939, 
        n14938, n14934, n14933, n14932, n14931, n14930, n14929, 
        n76_adj_5521, n79_adj_5522, n82_adj_5523, n85_adj_5524, n88_adj_5525, 
        n91_adj_5526, n94_adj_5527, n97_adj_5528, n100_adj_5529, n103_adj_5530, 
        n106_adj_5531, n109_adj_5532, n112_adj_5533, n115_adj_5534, 
        n118_adj_5535, n17027, n17293, n17635, n17573, n17572, n17098, 
        n45_adj_5536, n48_adj_5537, n51_adj_5538, n54_adj_5539, n57_adj_5540, 
        n60_adj_5541, n63_adj_5542, n66_adj_5543, n69_adj_5544, n72_adj_5545, 
        n75_adj_5546, n78_adj_5547, n81_adj_5548, n84_adj_5549, n87_adj_5550, 
        n90_adj_5551, n40, n49, n16740, n48_adj_5552, n51_adj_5553, 
        n54_adj_5554, n57_adj_5555, n60_adj_5556, n63_adj_5557, n66_adj_5558, 
        n69_adj_5559, n72_adj_5560, n75_adj_5561, n17317, n78_adj_5562, 
        n81_adj_5563, n84_adj_5564, n87_adj_5565, n90_adj_5566, n93_adj_5567, 
        n96_adj_5568, n99_adj_5569, n102_adj_5570, n105_adj_5571, n108_adj_5572, 
        n111_adj_5573, n114_adj_5574, n117_adj_5575, n120_adj_5576, 
        n123_adj_5577, n126_adj_5578, n129_adj_5579, n132_adj_5580, 
        n135_adj_5581, n138_adj_5582, n141_adj_5583, n144_adj_5584, 
        n147_adj_5585, n150_adj_5586, n153_adj_5587, n156_adj_5588, 
        n159_adj_5589, n162_adj_5590, n165_adj_5591, n168_adj_5592, 
        n171_adj_5593, n174_adj_5594, n177_adj_5595, n180_adj_5596, 
        n183_adj_5597, clk_80mhz_enable_1460, n17784, n14927, n124, 
        n14926, n127, n130_adj_5598, n133_adj_5599, n136_adj_5600, 
        n139_adj_5601, n142_adj_5602, n145_adj_5603, n148_adj_5604, 
        n151_adj_5605, n154_adj_5606, n14925, n157_adj_5607, n14924, 
        n160_adj_5608, n163_adj_5609, n166_adj_5610, n14923, n169_adj_5611, 
        n14922, n172_adj_5612, n14921, n175_adj_5613, n178_adj_5614, 
        n181_adj_5615, n16818, n184_adj_5616, n187_adj_5617, n190_adj_5618, 
        n193_adj_5619, n196_adj_5620, n199_adj_5621, n202_adj_5622, 
        n205_adj_5623, n208_adj_5624, n211_adj_5625, n214_adj_5626, 
        n217_adj_5627, n220_adj_5628, n223_adj_5629, n226_adj_5630, 
        n229_adj_5631, n232_adj_5632, n235_adj_5633, n238_adj_5634, 
        n241_adj_5635, n244_adj_5636, n247_adj_5637, n250_adj_5638, 
        n253_adj_5639, n256_adj_5640, n259_adj_5641, n262_adj_5642, 
        n265_adj_5643, n268_adj_5644, n271_adj_5645, n274_adj_5646, 
        n277_adj_5647, n280_adj_5648, n283_adj_5649, n286_adj_5650, 
        n289_adj_5651, n292_adj_5652, n295_adj_5653, n14920, n298_adj_5654, 
        n301_adj_5655, n14919, clk_80mhz_enable_45, n14918, n14917, 
        n17622, n14916, n17449, n17621, n17618, n17634, n16930, 
        n14915, n17648, n17647, n14914, n17646, n14913, n14912, 
        n14911, n14909, n12966, n17633, n17632, n13169, n17631, 
        n17522, n17521, cout_adj_5656, n14904, n14903, n14874, n14906, 
        n14907, n17630, n14899, n14902, n14901, n14900, n14910, 
        n14908, n17629, n14905;
    
    VHI i2 (.Z(VCC_net));
    CCU2C _add_1_1439_add_4_2 (.A0(d4_adj_5670[0]), .B0(d3_adj_5669[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[1]), .B1(d3_adj_5669[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15981), .S1(d4_71__N_634_adj_5686[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1439_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[36]), .B1(d7[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15921), .S1(n183_adj_4924));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1637_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_29 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15842), .COUT(n15843), .S0(n100), .S1(n97));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_29.INJECT1_1 = "NO";
    Mixer Mixer1 (.MixerOutSin({MixerOutSin}), .clk_80mhz(clk_80mhz), .DiffOut_c(DiffOut_c), 
          .MixerOutCos({MixerOutCos}), .RFIn_c(RFIn_c), .\LOCosine[3] (LOCosine[3]), 
          .MixerOutCos_11__N_250({MixerOutCos_11__N_250}), .\LOSine[1] (LOSine[1]), 
          .MixerOutSin_11__N_236({MixerOutSin_11__N_236}), .\LOCosine[1] (LOCosine[1]), 
          .\LOCosine[4] (LOCosine[4]), .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), 
          .\LOCosine[7] (LOCosine[7]), .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), 
          .\LOCosine[10] (LOCosine[10]), .\LOCosine[11] (LOCosine[11]), 
          .\LOCosine[12] (LOCosine[12]), .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), 
          .\LOSine[10] (LOSine[10]), .\LOSine[9] (LOSine[9]), .\LOSine[8] (LOSine[8]), 
          .\LOSine[7] (LOSine[7]), .\LOSine[6] (LOSine[6]), .\LOSine[5] (LOSine[5]), 
          .\LOSine[4] (LOSine[4]), .\LOSine[3] (LOSine[3]), .\LOSine[2] (LOSine[2]), 
          .\LOCosine[2] (LOCosine[2])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(166[7] 174[2])
    CCU2C _add_1_1484_add_4_27 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15841), .COUT(n15842), .S0(n106), .S1(n103));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_25 (.A0(d7_adj_5674[58]), .B0(cout_adj_5254), 
          .C0(n117_adj_5318), .D0(n15_adj_4641), .A1(d7_adj_5674[59]), 
          .B1(cout_adj_5254), .C1(n114_adj_5317), .D1(n14_adj_4642), .CIN(n16203), 
          .COUT(n16204), .S0(d8_71__N_1603_adj_5701[58]), .S1(d8_71__N_1603_adj_5701[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_3 (.A0(d6_adj_5672[36]), .B0(cout_adj_5179), 
          .C0(n183_adj_5304), .D0(n37_adj_4656), .A1(d6_adj_5672[37]), 
          .B1(cout_adj_5179), .C1(n180_adj_5303), .D1(n36_adj_4657), .CIN(n15961), 
          .COUT(n15962), .S0(d7_71__N_1531_adj_5700[36]), .S1(d7_71__N_1531_adj_5700[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15998), .S0(cout_adj_5136));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1439_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1439_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_34 (.A0(d4_adj_5670[32]), .B0(d3_adj_5669[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[33]), .B1(d3_adj_5669[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15996), .COUT(n15997), .S0(d4_71__N_634_adj_5686[32]), 
          .S1(d4_71__N_634_adj_5686[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_36 (.A0(d4_adj_5670[34]), .B0(d3_adj_5669[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[35]), .B1(d3_adj_5669[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15997), .COUT(n15998), .S0(d4_71__N_634_adj_5686[34]), 
          .S1(d4_71__N_634_adj_5686[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_36.INJECT1_1 = "NO";
    FD1S3AX o_Rx_DV_40 (.D(o_Rx_DV1), .CK(clk_80mhz), .Q(o_Rx_DV));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_DV_40.GSR = "ENABLED";
    CCU2C _add_1_1442_add_4_20 (.A0(d5_adj_5671[18]), .B0(d4_adj_5670[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[19]), .B1(d4_adj_5670[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15948), .COUT(n15949), .S0(d5_71__N_706_adj_5687[18]), 
          .S1(d5_71__N_706_adj_5687[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_20.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    CCU2C _add_1_1439_add_4_30 (.A0(d4_adj_5670[28]), .B0(d3_adj_5669[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[29]), .B1(d3_adj_5669[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15994), .COUT(n15995), .S0(d4_71__N_634_adj_5686[28]), 
          .S1(d4_71__N_634_adj_5686[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_30.INJECT1_1 = "NO";
    LUT4 mux_325_i21_4_lut (.A(n11953), .B(n259), .C(n17625), .D(n2571), 
         .Z(n2350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i21_4_lut.init = 16'hcfca;
    CCU2C _add_1_1484_add_4_25 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15840), .COUT(n15841), .S0(n112), .S1(n109));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_25.INJECT1_1 = "NO";
    PWM PWM1 (.\DataInReg[0] (DataInReg[0]), .clk_80mhz(clk_80mhz), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
        .counter({counter}), .\DemodOut[9] (DemodOut[9]), .\DataInReg[1] (DataInReg[1]), 
        .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg[2] (DataInReg[2]), 
        .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg[3] (DataInReg[3]), 
        .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg[4] (DataInReg[4]), 
        .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg[5] (DataInReg[5]), 
        .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg[6] (DataInReg[6]), 
        .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg[7] (DataInReg[7]), 
        .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg[8] (DataInReg[8]), 
        .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DataInReg[9] (DataInReg[9]), 
        .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(195[5] 201[2])
    CCU2C _add_1_1442_add_4_34 (.A0(d5_adj_5671[32]), .B0(d4_adj_5670[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[33]), .B1(d4_adj_5670[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15955), .COUT(n15956), .S0(d5_71__N_706_adj_5687[32]), 
          .S1(d5_71__N_706_adj_5687[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_23 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15839), .COUT(n15840), .S0(n118), .S1(n115));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_22 (.A0(d5_adj_5671[20]), .B0(d4_adj_5670[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[21]), .B1(d4_adj_5670[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15949), .COUT(n15950), .S0(d5_71__N_706_adj_5687[20]), 
          .S1(d5_71__N_706_adj_5687[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_21 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15838), .COUT(n15839));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_24 (.A0(d5_adj_5671[22]), .B0(d4_adj_5670[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[23]), .B1(d4_adj_5670[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15950), .COUT(n15951), .S0(d5_71__N_706_adj_5687[22]), 
          .S1(d5_71__N_706_adj_5687[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_19 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15837), .COUT(n15838));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_19.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_14 (.A0(MultResult2[12]), .B0(MultResult1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[13]), .B1(MultResult1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15800), .COUT(n15801), .S0(n90_adj_5166), 
          .S1(n87_adj_5165));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_14.INIT0 = 16'h666a;
    defparam ISquare_add_4_14.INIT1 = 16'h666a;
    defparam ISquare_add_4_14.INJECT1_0 = "NO";
    defparam ISquare_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_37 (.A0(d8_adj_5676[70]), .B0(cout_adj_5216), 
          .C0(n81), .D0(n3_adj_4615), .A1(d8_adj_5676[71]), .B1(cout_adj_5216), 
          .C1(n78), .D1(n2_adj_4616), .CIN(n15591), .S0(d9_71__N_1675_adj_5702[70]), 
          .S1(d9_71__N_1675_adj_5702[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_29 (.A0(d4_adj_5670[62]), .B0(cout_adj_5137), 
          .C0(n105), .D0(d5_adj_5671[62]), .A1(d4_adj_5670[63]), .B1(cout_adj_5137), 
          .C1(n102), .D1(d5_adj_5671[63]), .CIN(n15788), .COUT(n15789), 
          .S0(d5_71__N_706_adj_5687[62]), .S1(d5_71__N_706_adj_5687[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_26 (.A0(d5_adj_5671[24]), .B0(d4_adj_5670[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[25]), .B1(d4_adj_5670[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15951), .COUT(n15952), .S0(d5_71__N_706_adj_5687[24]), 
          .S1(d5_71__N_706_adj_5687[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_28 (.A0(d5_adj_5671[26]), .B0(d4_adj_5670[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[27]), .B1(d4_adj_5670[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15952), .COUT(n15953), .S0(d5_71__N_706_adj_5687[26]), 
          .S1(d5_71__N_706_adj_5687[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_17 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15836), .COUT(n15837));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_15 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15835), .COUT(n15836));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_35 (.A0(d8_adj_5676[68]), .B0(cout_adj_5216), 
          .C0(n87), .D0(n5_adj_4613), .A1(d8_adj_5676[69]), .B1(cout_adj_5216), 
          .C1(n84), .D1(n4_adj_4614), .CIN(n15590), .COUT(n15591), .S0(d9_71__N_1675_adj_5702[68]), 
          .S1(d9_71__N_1675_adj_5702[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_35.INJECT1_1 = "NO";
    FD1P3AX CICGain__i1 (.D(o_Rx_Byte[0]), .SP(clk_80mhz_enable_1408), .CK(clk_80mhz), 
            .Q(CICGain[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam CICGain__i1.GSR = "ENABLED";
    CCU2C _add_1_1475_add_4_23 (.A0(d7_adj_5674[56]), .B0(cout_adj_5254), 
          .C0(n123_adj_5320), .D0(n17_adj_4639), .A1(d7_adj_5674[57]), 
          .B1(cout_adj_5254), .C1(n120_adj_5319), .D1(n16_adj_4640), .CIN(n16202), 
          .COUT(n16203), .S0(d8_71__N_1603_adj_5701[56]), .S1(d8_71__N_1603_adj_5701[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_18 (.A0(d4_adj_5670[16]), .B0(d3_adj_5669[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[17]), .B1(d3_adj_5669[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15988), .COUT(n15989), .S0(d4_71__N_634_adj_5686[16]), 
          .S1(d4_71__N_634_adj_5686[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_18.INJECT1_1 = "NO";
    LUT4 mux_325_i22_4_lut (.A(n2549), .B(n256), .C(n17625), .D(n2571), 
         .Z(n2349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i22_4_lut.init = 16'hcfca;
    CCU2C _add_1_1439_add_4_32 (.A0(d4_adj_5670[30]), .B0(d3_adj_5669[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[31]), .B1(d3_adj_5669[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15995), .COUT(n15996), .S0(d4_71__N_634_adj_5686[30]), 
          .S1(d4_71__N_634_adj_5686[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_33 (.A0(d8_adj_5676[66]), .B0(cout_adj_5216), 
          .C0(n93_adj_4813), .D0(n7_adj_4611), .A1(d8_adj_5676[67]), .B1(cout_adj_5216), 
          .C1(n90), .D1(n6_adj_4612), .CIN(n15589), .COUT(n15590), .S0(d9_71__N_1675_adj_5702[66]), 
          .S1(d9_71__N_1675_adj_5702[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_21 (.A0(d7_adj_5674[54]), .B0(cout_adj_5254), 
          .C0(n129_adj_5322), .D0(n19_adj_4637), .A1(d7_adj_5674[55]), 
          .B1(cout_adj_5254), .C1(n126_adj_5321), .D1(n18_adj_4638), .CIN(n16201), 
          .COUT(n16202), .S0(d8_71__N_1603_adj_5701[54]), .S1(d8_71__N_1603_adj_5701[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15957), .S0(cout_adj_5137));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1442_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1442_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_16 (.A0(d4_adj_5670[14]), .B0(d3_adj_5669[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[15]), .B1(d3_adj_5669[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15987), .COUT(n15988), .S0(d4_71__N_634_adj_5686[14]), 
          .S1(d4_71__N_634_adj_5686[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_32 (.A0(d5_adj_5671[30]), .B0(d4_adj_5670[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[31]), .B1(d4_adj_5670[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15954), .COUT(n15955), .S0(d5_71__N_706_adj_5687[30]), 
          .S1(d5_71__N_706_adj_5687[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_14 (.A0(d4_adj_5670[12]), .B0(d3_adj_5669[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[13]), .B1(d3_adj_5669[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15986), .COUT(n15987), .S0(d4_71__N_634_adj_5686[12]), 
          .S1(d4_71__N_634_adj_5686[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_12 (.A0(d4_adj_5670[10]), .B0(d3_adj_5669[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[11]), .B1(d3_adj_5669[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15985), .COUT(n15986), .S0(d4_71__N_634_adj_5686[10]), 
          .S1(d4_71__N_634_adj_5686[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_10 (.A0(d4_adj_5670[8]), .B0(d3_adj_5669[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[9]), .B1(d3_adj_5669[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15984), .COUT(n15985), .S0(d4_71__N_634_adj_5686[8]), 
          .S1(d4_71__N_634_adj_5686[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_13 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15834), .COUT(n15835));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_8 (.A0(d4_adj_5670[6]), .B0(d3_adj_5669[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[7]), .B1(d3_adj_5669[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15983), .COUT(n15984), .S0(d4_71__N_634_adj_5686[6]), 
          .S1(d4_71__N_634_adj_5686[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_27 (.A0(d4_adj_5670[60]), .B0(cout_adj_5137), 
          .C0(n111), .D0(d5_adj_5671[60]), .A1(d4_adj_5670[61]), .B1(cout_adj_5137), 
          .C1(n108), .D1(d5_adj_5671[61]), .CIN(n15787), .COUT(n15788), 
          .S0(d5_71__N_706_adj_5687[60]), .S1(d5_71__N_706_adj_5687[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_37 (.A0(d7[70]), .B0(cout_adj_5088), .C0(n81_adj_4890), 
          .D0(n3_adj_4692), .A1(d7[71]), .B1(cout_adj_5088), .C1(n78_adj_4889), 
          .D1(n2_adj_4693), .CIN(n15919), .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_16 (.A0(d5_adj_5671[14]), .B0(d4_adj_5670[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[15]), .B1(d4_adj_5670[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15946), .COUT(n15947), .S0(d5_71__N_706_adj_5687[14]), 
          .S1(d5_71__N_706_adj_5687[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_11 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15833), .COUT(n15834));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_9 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15832), .COUT(n15833));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_7 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15831), .COUT(n15832));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_5 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15830), .COUT(n15831));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_31 (.A0(d8_adj_5676[64]), .B0(cout_adj_5216), 
          .C0(n99_adj_4789), .D0(n9_adj_4609), .A1(d8_adj_5676[65]), .B1(cout_adj_5216), 
          .C1(n96_adj_4790), .D1(n8_adj_4610), .CIN(n15588), .COUT(n15589), 
          .S0(d9_71__N_1675_adj_5702[64]), .S1(d9_71__N_1675_adj_5702[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5179), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15961));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1478_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1478_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_6 (.A0(d4_adj_5670[4]), .B0(d3_adj_5669[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[5]), .B1(d3_adj_5669[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15982), .COUT(n15983), .S0(d4_71__N_634_adj_5686[4]), 
          .S1(d4_71__N_634_adj_5686[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_3 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15829), .COUT(n15830));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_29 (.A0(d8_adj_5676[62]), .B0(cout_adj_5216), 
          .C0(n105_adj_4787), .D0(n11_adj_4607), .A1(d8_adj_5676[63]), 
          .B1(cout_adj_5216), .C1(n102_adj_4788), .D1(n10_adj_4608), .CIN(n15587), 
          .COUT(n15588), .S0(d9_71__N_1675_adj_5702[62]), .S1(d9_71__N_1675_adj_5702[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_4 (.A0(d4_adj_5670[2]), .B0(d3_adj_5669[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[3]), .B1(d3_adj_5669[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15981), .COUT(n15982), .S0(d4_71__N_634_adj_5686[2]), 
          .S1(d4_71__N_634_adj_5686[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_19 (.A0(d7_adj_5674[52]), .B0(cout_adj_5254), 
          .C0(n135_adj_5324), .D0(n21_adj_4635), .A1(d7_adj_5674[53]), 
          .B1(cout_adj_5254), .C1(n132_adj_5323), .D1(n20_adj_4636), .CIN(n16200), 
          .COUT(n16201), .S0(d8_71__N_1603_adj_5701[52]), .S1(d8_71__N_1603_adj_5701[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_17 (.A0(d7_adj_5674[50]), .B0(cout_adj_5254), 
          .C0(n141_adj_5326), .D0(n23_adj_4633), .A1(d7_adj_5674[51]), 
          .B1(cout_adj_5254), .C1(n138_adj_5325), .D1(n22_adj_4634), .CIN(n16199), 
          .COUT(n16200), .S0(d8_71__N_1603_adj_5701[50]), .S1(d8_71__N_1603_adj_5701[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_15 (.A0(d7_adj_5674[48]), .B0(cout_adj_5254), 
          .C0(n147_adj_5328), .D0(n25_adj_4631), .A1(d7_adj_5674[49]), 
          .B1(cout_adj_5254), .C1(n144_adj_5327), .D1(n24_adj_4632), .CIN(n16198), 
          .COUT(n16199), .S0(d8_71__N_1603_adj_5701[48]), .S1(d8_71__N_1603_adj_5701[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_13 (.A0(d7_adj_5674[46]), .B0(cout_adj_5254), 
          .C0(n153_adj_5330), .D0(n27_adj_4629), .A1(d7_adj_5674[47]), 
          .B1(cout_adj_5254), .C1(n150_adj_5329), .D1(n26_adj_4630), .CIN(n16197), 
          .COUT(n16198), .S0(d8_71__N_1603_adj_5701[46]), .S1(d8_71__N_1603_adj_5701[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_11 (.A0(d7_adj_5674[44]), .B0(cout_adj_5254), 
          .C0(n159_adj_5332), .D0(n29_adj_4627), .A1(d7_adj_5674[45]), 
          .B1(cout_adj_5254), .C1(n156_adj_5331), .D1(n28_adj_4628), .CIN(n16196), 
          .COUT(n16197), .S0(d8_71__N_1603_adj_5701[44]), .S1(d8_71__N_1603_adj_5701[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_9 (.A0(d7_adj_5674[42]), .B0(cout_adj_5254), 
          .C0(n165_adj_5334), .D0(n31_adj_4624), .A1(d7_adj_5674[43]), 
          .B1(cout_adj_5254), .C1(n162_adj_5333), .D1(n30_adj_4626), .CIN(n16195), 
          .COUT(n16196), .S0(d8_71__N_1603_adj_5701[42]), .S1(d8_71__N_1603_adj_5701[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_7 (.A0(d7_adj_5674[40]), .B0(cout_adj_5254), 
          .C0(n171_adj_5336), .D0(n33_adj_4622), .A1(d7_adj_5674[41]), 
          .B1(cout_adj_5254), .C1(n168_adj_5335), .D1(n32_adj_4623), .CIN(n16194), 
          .COUT(n16195), .S0(d8_71__N_1603_adj_5701[40]), .S1(d8_71__N_1603_adj_5701[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_5 (.A0(d7_adj_5674[38]), .B0(cout_adj_5254), 
          .C0(n177_adj_5338), .D0(n35_adj_4620), .A1(d7_adj_5674[39]), 
          .B1(cout_adj_5254), .C1(n174_adj_5337), .D1(n34_adj_4621), .CIN(n16193), 
          .COUT(n16194), .S0(d8_71__N_1603_adj_5701[38]), .S1(d8_71__N_1603_adj_5701[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_3 (.A0(d7_adj_5674[36]), .B0(cout_adj_5254), 
          .C0(n183_adj_5340), .D0(n37_adj_4618), .A1(d7_adj_5674[37]), 
          .B1(cout_adj_5254), .C1(n180_adj_5339), .D1(n36_adj_4619), .CIN(n16192), 
          .COUT(n16193), .S0(d8_71__N_1603_adj_5701[36]), .S1(d8_71__N_1603_adj_5701[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5254), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16192));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1475_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1475_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_29 (.A0(d6_adj_5672[62]), .B0(cout_adj_5179), 
          .C0(n105_adj_5278), .D0(n11_adj_4684), .A1(d6_adj_5672[63]), 
          .B1(cout_adj_5179), .C1(n102_adj_5277), .D1(n10_adj_4683), .CIN(n15974), 
          .COUT(n15975), .S0(d7_71__N_1531_adj_5700[62]), .S1(d7_71__N_1531_adj_5700[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15829));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1484_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_1.INJECT1_1 = "NO";
    LUT4 i5098_2_lut_rep_173 (.A(ISquare[23]), .B(ISquare[22]), .Z(n17642)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam i5098_2_lut_rep_173.init = 16'heeee;
    LUT4 i5142_1_lut_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n40)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam i5142_1_lut_2_lut_3_lut.init = 16'h0101;
    CCU2C _add_1_1472_add_4_27 (.A0(d8_adj_5676[60]), .B0(cout_adj_5216), 
          .C0(n111_adj_4785), .D0(n13_adj_4605), .A1(d8_adj_5676[61]), 
          .B1(cout_adj_5216), .C1(n108_adj_4786), .D1(n12_adj_4606), .CIN(n15586), 
          .COUT(n15587), .S0(d9_71__N_1675_adj_5702[60]), .S1(d9_71__N_1675_adj_5702[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_27.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_166_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n17635)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam i1_2_lut_rep_166_3_lut.init = 16'hfefe;
    CCU2C _add_1_1466_add_4_35 (.A0(d7[68]), .B0(cout_adj_5088), .C0(n87_adj_4892), 
          .D0(n5_adj_4690), .A1(d7[69]), .B1(cout_adj_5088), .C1(n84_adj_4891), 
          .D1(n4_adj_4691), .CIN(n15918), .COUT(n15919), .S0(d8_71__N_1603[68]), 
          .S1(d8_71__N_1603[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_19 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n135_adj_5109), .D0(d1[52]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n132_adj_5108), .D1(d1[53]), .CIN(n15858), .COUT(n15859), 
          .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_33 (.A0(d7[66]), .B0(cout_adj_5088), .C0(n93_adj_4894), 
          .D0(n7_adj_4687), .A1(d7[67]), .B1(cout_adj_5088), .C1(n90_adj_4893), 
          .D1(n6_adj_4689), .CIN(n15917), .COUT(n15918), .S0(d8_71__N_1603[66]), 
          .S1(d8_71__N_1603[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_17 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n141_adj_5111), .D0(d1[50]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n138_adj_5110), .D1(d1[51]), .CIN(n15857), .COUT(n15858), 
          .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_12 (.A0(d5_adj_5671[10]), .B0(d4_adj_5670[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[11]), .B1(d4_adj_5670[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15944), .COUT(n15945), .S0(d5_71__N_706_adj_5687[10]), 
          .S1(d5_71__N_706_adj_5687[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_37 (.A0(d8[70]), .B0(cout_adj_5000), .C0(n81_adj_5002), 
          .D0(n3_adj_4834), .A1(d8[71]), .B1(cout_adj_5000), .C1(n78_adj_5001), 
          .D1(n2_adj_4835), .CIN(n15827), .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_10 (.A0(d5_adj_5671[8]), .B0(d4_adj_5670[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[9]), .B1(d4_adj_5670[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15943), .COUT(n15944), .S0(d5_71__N_706_adj_5687[8]), 
          .S1(d5_71__N_706_adj_5687[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_4 (.A0(d5_adj_5671[2]), .B0(d4_adj_5670[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[3]), .B1(d4_adj_5670[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15940), .COUT(n15941), .S0(d5_71__N_706_adj_5687[2]), 
          .S1(d5_71__N_706_adj_5687[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_38 (.A0(d_d7[71]), .B0(d7[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15938), .S0(n78_adj_4889));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1637_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_31 (.A0(d7[64]), .B0(cout_adj_5088), .C0(n99_adj_4896), 
          .D0(n9_adj_4655), .A1(d7[65]), .B1(cout_adj_5088), .C1(n96_adj_4895), 
          .D1(n8_adj_4658), .CIN(n15916), .COUT(n15917), .S0(d8_71__N_1603[64]), 
          .S1(d8_71__N_1603[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_2 (.A0(d5_adj_5671[0]), .B0(d4_adj_5670[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[1]), .B1(d4_adj_5670[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15940), .S1(d5_71__N_706_adj_5687[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1442_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_8 (.A0(d5_adj_5671[6]), .B0(d4_adj_5670[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[7]), .B1(d4_adj_5670[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15942), .COUT(n15943), .S0(d5_71__N_706_adj_5687[6]), 
          .S1(d5_71__N_706_adj_5687[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_36 (.A0(d_d7[69]), .B0(d7[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[70]), .B1(d7[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15937), .COUT(n15938), .S0(n84_adj_4891), .S1(n81_adj_4890));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_6 (.A0(d5_adj_5671[4]), .B0(d4_adj_5670[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[5]), .B1(d4_adj_5670[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15941), .COUT(n15942), .S0(d5_71__N_706_adj_5687[4]), 
          .S1(d5_71__N_706_adj_5687[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_25 (.A0(d8_adj_5676[58]), .B0(cout_adj_5216), 
          .C0(n117_adj_4783), .D0(n15_adj_4603), .A1(d8_adj_5676[59]), 
          .B1(cout_adj_5216), .C1(n114_adj_4784), .D1(n14_adj_4604), .CIN(n15585), 
          .COUT(n15586), .S0(d9_71__N_1675_adj_5702[58]), .S1(d9_71__N_1675_adj_5702[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_23 (.A0(d8_adj_5676[56]), .B0(cout_adj_5216), 
          .C0(n123_adj_4767), .D0(n17_adj_4601), .A1(d8_adj_5676[57]), 
          .B1(cout_adj_5216), .C1(n120_adj_4782), .D1(n16_adj_4602), .CIN(n15584), 
          .COUT(n15585), .S0(d9_71__N_1675_adj_5702[56]), .S1(d9_71__N_1675_adj_5702[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_21 (.A0(d8_adj_5676[54]), .B0(cout_adj_5216), 
          .C0(n129_adj_4765), .D0(n19_adj_4599), .A1(d8_adj_5676[55]), 
          .B1(cout_adj_5216), .C1(n126_adj_4766), .D1(n18_adj_4600), .CIN(n15583), 
          .COUT(n15584), .S0(d9_71__N_1675_adj_5702[54]), .S1(d9_71__N_1675_adj_5702[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_29 (.A0(d7[62]), .B0(cout_adj_5088), .C0(n105_adj_4898), 
          .D0(n11_adj_4617), .A1(d7[63]), .B1(cout_adj_5088), .C1(n102_adj_4897), 
          .D1(n10_adj_4625), .CIN(n15915), .COUT(n15916), .S0(d8_71__N_1603[62]), 
          .S1(d8_71__N_1603[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_19 (.A0(d8_adj_5676[52]), .B0(cout_adj_5216), 
          .C0(n135_adj_4749), .D0(n21_adj_4597), .A1(d8_adj_5676[53]), 
          .B1(cout_adj_5216), .C1(n132_adj_4750), .D1(n20_adj_4598), .CIN(n15582), 
          .COUT(n15583), .S0(d9_71__N_1675_adj_5702[52]), .S1(d9_71__N_1675_adj_5702[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_17 (.A0(d8_adj_5676[50]), .B0(cout_adj_5216), 
          .C0(n141_adj_4747), .D0(n23_adj_4595), .A1(d8_adj_5676[51]), 
          .B1(cout_adj_5216), .C1(n138_adj_4748), .D1(n22_adj_4596), .CIN(n15581), 
          .COUT(n15582), .S0(d9_71__N_1675_adj_5702[50]), .S1(d9_71__N_1675_adj_5702[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_25 (.A0(d4_adj_5670[58]), .B0(cout_adj_5137), 
          .C0(n117), .D0(d5_adj_5671[58]), .A1(d4_adj_5670[59]), .B1(cout_adj_5137), 
          .C1(n114), .D1(d5_adj_5671[59]), .CIN(n15786), .COUT(n15787), 
          .S0(d5_71__N_706_adj_5687[58]), .S1(d5_71__N_706_adj_5687[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_27 (.A0(d7[60]), .B0(cout_adj_5088), .C0(n111_adj_4900), 
          .D0(n13_adj_4579), .A1(d7[61]), .B1(cout_adj_5088), .C1(n108_adj_4899), 
          .D1(n12_adj_4592), .CIN(n15914), .COUT(n15915), .S0(d8_71__N_1603[60]), 
          .S1(d8_71__N_1603[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_27.INJECT1_1 = "NO";
    LUT4 i5126_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n14874)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam i5126_2_lut_3_lut.init = 16'h0e0e;
    CCU2C _add_1_1478_add_4_37 (.A0(d6_adj_5672[70]), .B0(cout_adj_5179), 
          .C0(n81_adj_5270), .D0(n3), .A1(d6_adj_5672[71]), .B1(cout_adj_5179), 
          .C1(n78_adj_5269), .D1(n2), .CIN(n15978), .S0(d7_71__N_1531_adj_5700[70]), 
          .S1(d7_71__N_1531_adj_5700[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_25 (.A0(d7[58]), .B0(cout_adj_5088), .C0(n117_adj_4902), 
          .D0(n15_adj_4577), .A1(d7[59]), .B1(cout_adj_5088), .C1(n114_adj_4901), 
          .D1(n14_adj_4578), .CIN(n15913), .COUT(n15914), .S0(d8_71__N_1603[58]), 
          .S1(d8_71__N_1603[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_15 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n147_adj_5113), .D0(d1[48]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n144_adj_5112), .D1(d1[49]), .CIN(n15856), .COUT(n15857), 
          .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_34 (.A0(d_d7[67]), .B0(d7[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[68]), .B1(d7[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15936), .COUT(n15937), .S0(n90_adj_4893), .S1(n87_adj_4892));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_32 (.A0(d_d7[65]), .B0(d7[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[66]), .B1(d7[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15935), .COUT(n15936), .S0(n96_adj_4895), .S1(n93_adj_4894));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_30 (.A0(d_d7[63]), .B0(d7[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[64]), .B1(d7[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15934), .COUT(n15935), .S0(n102_adj_4897), .S1(n99_adj_4896));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_13 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n153_adj_5115), .D0(d1[46]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n150_adj_5114), .D1(d1[47]), .CIN(n15855), .COUT(n15856), 
          .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_13.INJECT1_1 = "NO";
    LUT4 i5116_1_lut_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n49)) /* synthesis lut_function=(!(A+(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam i5116_1_lut_2_lut.init = 16'h1111;
    CCU2C _add_1_1637_add_4_28 (.A0(d_d7[61]), .B0(d7[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[62]), .B1(d7[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15933), .COUT(n15934), .S0(n108_adj_4899), .S1(n105_adj_4898));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_24 (.A0(d_d7[57]), .B0(d7[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[58]), .B1(d7[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15931), .COUT(n15932), .S0(n120_adj_4903), .S1(n117_adj_4902));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_26 (.A0(d_d7[59]), .B0(d7[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[60]), .B1(d7[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15932), .COUT(n15933), .S0(n114_adj_4901), .S1(n111_adj_4900));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_23 (.A0(d7[56]), .B0(cout_adj_5088), .C0(n123_adj_4904), 
          .D0(n17_adj_4575), .A1(d7[57]), .B1(cout_adj_5088), .C1(n120_adj_4903), 
          .D1(n16_adj_4576), .CIN(n15912), .COUT(n15913), .S0(d8_71__N_1603[56]), 
          .S1(d8_71__N_1603[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_23.INJECT1_1 = "NO";
    LUT4 i359_2_lut_3_lut_4_lut_4_lut (.A(n17751), .B(n17634), .C(o_Rx_Byte[4]), 
         .D(o_Rx_Byte[0]), .Z(n2571)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i359_2_lut_3_lut_4_lut_4_lut.init = 16'h0400;
    CCU2C _add_1_1472_add_4_15 (.A0(d8_adj_5676[48]), .B0(cout_adj_5216), 
          .C0(n147_adj_4745), .D0(n25_adj_4593), .A1(d8_adj_5676[49]), 
          .B1(cout_adj_5216), .C1(n144_adj_4746), .D1(n24_adj_4594), .CIN(n15580), 
          .COUT(n15581), .S0(d9_71__N_1675_adj_5702[48]), .S1(d9_71__N_1675_adj_5702[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_35 (.A0(d6_adj_5672[68]), .B0(cout_adj_5179), 
          .C0(n87_adj_5272), .D0(n5), .A1(d6_adj_5672[69]), .B1(cout_adj_5179), 
          .C1(n84_adj_5271), .D1(n4), .CIN(n15977), .COUT(n15978), .S0(d7_71__N_1531_adj_5700[68]), 
          .S1(d7_71__N_1531_adj_5700[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_13 (.A0(d8_adj_5676[46]), .B0(cout_adj_5216), 
          .C0(n153_adj_4743), .D0(n27_adj_4590), .A1(d8_adj_5676[47]), 
          .B1(cout_adj_5216), .C1(n150_adj_4744), .D1(n26_adj_4591), .CIN(n15579), 
          .COUT(n15580), .S0(d9_71__N_1675_adj_5702[46]), .S1(d9_71__N_1675_adj_5702[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_7 (.A0(d6_adj_5672[40]), .B0(cout_adj_5179), 
          .C0(n171_adj_5300), .D0(n33_adj_4661), .A1(d6_adj_5672[41]), 
          .B1(cout_adj_5179), .C1(n168_adj_5299), .D1(n32_adj_4662), .CIN(n15963), 
          .COUT(n15964), .S0(d7_71__N_1531_adj_5700[40]), .S1(d7_71__N_1531_adj_5700[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_7.INJECT1_1 = "NO";
    LUT4 CIC_out_clkSin_c_bdd_2_lut_6211_2_lut (.A(o_Rx_Byte[3]), .B(n17572), 
         .Z(n17573)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam CIC_out_clkSin_c_bdd_2_lut_6211_2_lut.init = 16'h4444;
    CCU2C _add_1_1478_add_4_33 (.A0(d6_adj_5672[66]), .B0(cout_adj_5179), 
          .C0(n93_adj_5274), .D0(n7), .A1(d6_adj_5672[67]), .B1(cout_adj_5179), 
          .C1(n90_adj_5273), .D1(n6), .CIN(n15976), .COUT(n15977), .S0(d7_71__N_1531_adj_5700[66]), 
          .S1(d7_71__N_1531_adj_5700[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_35 (.A0(d8[68]), .B0(cout_adj_5000), .C0(n87_adj_5004), 
          .D0(n5_adj_4832), .A1(d8[69]), .B1(cout_adj_5000), .C1(n84_adj_5003), 
          .D1(n4_adj_4833), .CIN(n15826), .COUT(n15827), .S0(d9_71__N_1675[68]), 
          .S1(d9_71__N_1675[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_33 (.A0(d8[66]), .B0(cout_adj_5000), .C0(n93_adj_5006), 
          .D0(n7_adj_4830), .A1(d8[67]), .B1(cout_adj_5000), .C1(n90_adj_5005), 
          .D1(n6_adj_4831), .CIN(n15825), .COUT(n15826), .S0(d9_71__N_1675[66]), 
          .S1(d9_71__N_1675[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_31 (.A0(d8[64]), .B0(cout_adj_5000), .C0(n99_adj_5008), 
          .D0(n9_adj_4828), .A1(d8[65]), .B1(cout_adj_5000), .C1(n96_adj_5007), 
          .D1(n8_adj_4829), .CIN(n15824), .COUT(n15825), .S0(d9_71__N_1675[64]), 
          .S1(d9_71__N_1675[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_11 (.A0(d8_adj_5676[44]), .B0(cout_adj_5216), 
          .C0(n159_adj_4741), .D0(n29_adj_4588), .A1(d8_adj_5676[45]), 
          .B1(cout_adj_5216), .C1(n156_adj_4742), .D1(n28_adj_4589), .CIN(n15578), 
          .COUT(n15579), .S0(d9_71__N_1675_adj_5702[44]), .S1(d9_71__N_1675_adj_5702[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_29 (.A0(d8[62]), .B0(cout_adj_5000), .C0(n105_adj_5010), 
          .D0(n11_adj_4826), .A1(d8[63]), .B1(cout_adj_5000), .C1(n102_adj_5009), 
          .D1(n10_adj_4827), .CIN(n15823), .COUT(n15824), .S0(d9_71__N_1675[62]), 
          .S1(d9_71__N_1675[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_9 (.A0(d8_adj_5676[42]), .B0(cout_adj_5216), 
          .C0(n165_adj_4739), .D0(n31_adj_4586), .A1(d8_adj_5676[43]), 
          .B1(cout_adj_5216), .C1(n162_adj_4740), .D1(n30_adj_4587), .CIN(n15577), 
          .COUT(n15578), .S0(d9_71__N_1675_adj_5702[42]), .S1(d9_71__N_1675_adj_5702[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_27 (.A0(d8[60]), .B0(cout_adj_5000), .C0(n111_adj_5012), 
          .D0(n13_adj_4824), .A1(d8[61]), .B1(cout_adj_5000), .C1(n108_adj_5011), 
          .D1(n12_adj_4825), .CIN(n15822), .COUT(n15823), .S0(d9_71__N_1675[60]), 
          .S1(d9_71__N_1675[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_31 (.A0(d6_adj_5672[64]), .B0(cout_adj_5179), 
          .C0(n99_adj_5276), .D0(n9_adj_4682), .A1(d6_adj_5672[65]), .B1(cout_adj_5179), 
          .C1(n96_adj_5275), .D1(n8_adj_4686), .CIN(n15975), .COUT(n15976), 
          .S0(d7_71__N_1531_adj_5700[64]), .S1(d7_71__N_1531_adj_5700[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_25 (.A0(d8[58]), .B0(cout_adj_5000), .C0(n117_adj_5014), 
          .D0(n15_adj_4822), .A1(d8[59]), .B1(cout_adj_5000), .C1(n114_adj_5013), 
          .D1(n14_adj_4823), .CIN(n15821), .COUT(n15822), .S0(d9_71__N_1675[58]), 
          .S1(d9_71__N_1675[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_23 (.A0(d8[56]), .B0(cout_adj_5000), .C0(n123_adj_5016), 
          .D0(n17_adj_4820), .A1(d8[57]), .B1(cout_adj_5000), .C1(n120_adj_5015), 
          .D1(n16_adj_4821), .CIN(n15820), .COUT(n15821), .S0(d9_71__N_1675[56]), 
          .S1(d9_71__N_1675[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_21 (.A0(d8[54]), .B0(cout_adj_5000), .C0(n129_adj_5018), 
          .D0(n19_adj_4818), .A1(d8[55]), .B1(cout_adj_5000), .C1(n126_adj_5017), 
          .D1(n18_adj_4819), .CIN(n15819), .COUT(n15820), .S0(d9_71__N_1675[54]), 
          .S1(d9_71__N_1675[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_19 (.A0(d8[52]), .B0(cout_adj_5000), .C0(n135_adj_5020), 
          .D0(n21_adj_4816), .A1(d8[53]), .B1(cout_adj_5000), .C1(n132_adj_5019), 
          .D1(n20_adj_4817), .CIN(n15818), .COUT(n15819), .S0(d9_71__N_1675[52]), 
          .S1(d9_71__N_1675[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_17 (.A0(d8[50]), .B0(cout_adj_5000), .C0(n141_adj_5022), 
          .D0(n23_adj_4814), .A1(d8[51]), .B1(cout_adj_5000), .C1(n138_adj_5021), 
          .D1(n22_adj_4815), .CIN(n15817), .COUT(n15818), .S0(d9_71__N_1675[50]), 
          .S1(d9_71__N_1675[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_15 (.A0(d8[48]), .B0(cout_adj_5000), .C0(n147_adj_5024), 
          .D0(n25_adj_4780), .A1(d8[49]), .B1(cout_adj_5000), .C1(n144_adj_5023), 
          .D1(n24_adj_4781), .CIN(n15816), .COUT(n15817), .S0(d9_71__N_1675[48]), 
          .S1(d9_71__N_1675[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_7 (.A0(d8_adj_5676[40]), .B0(cout_adj_5216), 
          .C0(n171_adj_4737), .D0(n33_adj_4584), .A1(d8_adj_5676[41]), 
          .B1(cout_adj_5216), .C1(n168_adj_4738), .D1(n32_adj_4585), .CIN(n15576), 
          .COUT(n15577), .S0(d9_71__N_1675_adj_5702[40]), .S1(d9_71__N_1675_adj_5702[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4999), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15850));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1448_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1448_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_13 (.A0(d8[46]), .B0(cout_adj_5000), .C0(n153_adj_5026), 
          .D0(n27_adj_4778), .A1(d8[47]), .B1(cout_adj_5000), .C1(n150_adj_5025), 
          .D1(n26_adj_4779), .CIN(n15815), .COUT(n15816), .S0(d9_71__N_1675[46]), 
          .S1(d9_71__N_1675[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_11 (.A0(d8[44]), .B0(cout_adj_5000), .C0(n159_adj_5028), 
          .D0(n29_adj_4776), .A1(d8[45]), .B1(cout_adj_5000), .C1(n156_adj_5027), 
          .D1(n28_adj_4777), .CIN(n15814), .COUT(n15815), .S0(d9_71__N_1675[44]), 
          .S1(d9_71__N_1675[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_9 (.A0(d8[42]), .B0(cout_adj_5000), .C0(n165_adj_5030), 
          .D0(n31_adj_4774), .A1(d8[43]), .B1(cout_adj_5000), .C1(n162_adj_5029), 
          .D1(n30_adj_4775), .CIN(n15813), .COUT(n15814), .S0(d9_71__N_1675[42]), 
          .S1(d9_71__N_1675[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_7 (.A0(d8[40]), .B0(cout_adj_5000), .C0(n171_adj_5032), 
          .D0(n33_adj_4772), .A1(d8[41]), .B1(cout_adj_5000), .C1(n168_adj_5031), 
          .D1(n32_adj_4773), .CIN(n15812), .COUT(n15813), .S0(d9_71__N_1675[40]), 
          .S1(d9_71__N_1675[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_5 (.A0(d8[38]), .B0(cout_adj_5000), .C0(n177_adj_5034), 
          .D0(n35_adj_4770), .A1(d8[39]), .B1(cout_adj_5000), .C1(n174_adj_5033), 
          .D1(n34_adj_4771), .CIN(n15811), .COUT(n15812), .S0(d9_71__N_1675[38]), 
          .S1(d9_71__N_1675[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_3 (.A0(d8[36]), .B0(cout_adj_5000), .C0(n183_adj_5036), 
          .D0(n37_adj_4768), .A1(d8[37]), .B1(cout_adj_5000), .C1(n180_adj_5035), 
          .D1(n36_adj_4769), .CIN(n15810), .COUT(n15811), .S0(d9_71__N_1675[36]), 
          .S1(d9_71__N_1675[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1487_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1487_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5000), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15810));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1487_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1487_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1487_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_1.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_26 (.A0(MultResult2[23]), .B0(MultResult1[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15806), .S0(n54_adj_5154));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_26.INIT0 = 16'h666a;
    defparam ISquare_add_4_26.INIT1 = 16'h0000;
    defparam ISquare_add_4_26.INJECT1_0 = "NO";
    defparam ISquare_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_5 (.A0(d8_adj_5676[38]), .B0(cout_adj_5216), 
          .C0(n177_adj_4735), .D0(n35_adj_4582), .A1(d8_adj_5676[39]), 
          .B1(cout_adj_5216), .C1(n174_adj_4736), .D1(n34_adj_4583), .CIN(n15575), 
          .COUT(n15576), .S0(d9_71__N_1675_adj_5702[38]), .S1(d9_71__N_1675_adj_5702[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_5.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_24 (.A0(MultResult2[22]), .B0(MultResult1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[23]), .B1(MultResult1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15805), .COUT(n15806), .S0(n60_adj_5156), 
          .S1(n57_adj_5155));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_24.INIT0 = 16'h666a;
    defparam ISquare_add_4_24.INIT1 = 16'h666a;
    defparam ISquare_add_4_24.INJECT1_0 = "NO";
    defparam ISquare_add_4_24.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_22 (.A0(MultResult2[20]), .B0(MultResult1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[21]), .B1(MultResult1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15804), .COUT(n15805), .S0(n66_adj_5158), 
          .S1(n63_adj_5157));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_22.INIT0 = 16'h666a;
    defparam ISquare_add_4_22.INIT1 = 16'h666a;
    defparam ISquare_add_4_22.INJECT1_0 = "NO";
    defparam ISquare_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_38 (.A0(d_d6_adj_5673[71]), .B0(d6_adj_5672[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16188), .S0(n78_adj_5269));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1625_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_22 (.A0(d_d7[55]), .B0(d7[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[56]), .B1(d7[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15930), .COUT(n15931), .S0(n126_adj_4905), .S1(n123_adj_4904));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_21 (.A0(d7[54]), .B0(cout_adj_5088), .C0(n129_adj_4906), 
          .D0(n19_adj_4573), .A1(d7[55]), .B1(cout_adj_5088), .C1(n126_adj_4905), 
          .D1(n18_adj_4574), .CIN(n15911), .COUT(n15912), .S0(d8_71__N_1603[54]), 
          .S1(d8_71__N_1603[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_14 (.A0(d_d7[47]), .B0(d7[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[48]), .B1(d7[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15926), .COUT(n15927), .S0(n150_adj_4913), .S1(n147_adj_4912));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_23 (.A0(d4_adj_5670[56]), .B0(cout_adj_5137), 
          .C0(n123), .D0(d5_adj_5671[56]), .A1(d4_adj_5670[57]), .B1(cout_adj_5137), 
          .C1(n120), .D1(d5_adj_5671[57]), .CIN(n15785), .COUT(n15786), 
          .S0(d5_71__N_706_adj_5687[56]), .S1(d5_71__N_706_adj_5687[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_23.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_12 (.A0(MultResult2[10]), .B0(MultResult1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[11]), .B1(MultResult1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15799), .COUT(n15800), .S0(n96_adj_5168), 
          .S1(n93_adj_5167));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_12.INIT0 = 16'h666a;
    defparam ISquare_add_4_12.INIT1 = 16'h666a;
    defparam ISquare_add_4_12.INJECT1_0 = "NO";
    defparam ISquare_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_3 (.A0(d8_adj_5676[36]), .B0(cout_adj_5216), 
          .C0(n183_adj_4733), .D0(n37_adj_4580), .A1(d8_adj_5676[37]), 
          .B1(cout_adj_5216), .C1(n180_adj_4734), .D1(n36_adj_4581), .CIN(n15574), 
          .COUT(n15575), .S0(d9_71__N_1675_adj_5702[36]), .S1(d9_71__N_1675_adj_5702[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1472_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1472_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_12 (.A0(d_d7[45]), .B0(d7[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[46]), .B1(d7[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15925), .COUT(n15926), .S0(n156_adj_4915), .S1(n153_adj_4914));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_3 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n183_adj_5125), .D0(d1[36]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n180_adj_5124), .D1(d1[37]), .CIN(n15850), .COUT(n15851), 
          .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_10 (.A0(d_d7[43]), .B0(d7[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[44]), .B1(d7[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15924), .COUT(n15925), .S0(n162_adj_4917), .S1(n159_adj_4916));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_20 (.A0(d_d7[53]), .B0(d7[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[54]), .B1(d7[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15929), .COUT(n15930), .S0(n132_adj_4907), .S1(n129_adj_4906));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_8 (.A0(d_d7[41]), .B0(d7[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[42]), .B1(d7[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15923), .COUT(n15924), .S0(n168_adj_4919), .S1(n165_adj_4918));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_27 (.A0(d6_adj_5672[60]), .B0(cout_adj_5179), 
          .C0(n111_adj_5280), .D0(n13_adj_4681), .A1(d6_adj_5672[61]), 
          .B1(cout_adj_5179), .C1(n108_adj_5279), .D1(n12_adj_4685), .CIN(n15973), 
          .COUT(n15974), .S0(d7_71__N_1531_adj_5700[60]), .S1(d7_71__N_1531_adj_5700[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_5 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n177_adj_5123), .D0(d1[38]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n174_adj_5122), .D1(d1[39]), .CIN(n15851), .COUT(n15852), 
          .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_11 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n159_adj_5117), .D0(d1[44]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n156_adj_5116), .D1(d1[45]), .CIN(n15854), .COUT(n15855), 
          .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_25 (.A0(d6_adj_5672[58]), .B0(cout_adj_5179), 
          .C0(n117_adj_5282), .D0(n15_adj_4679), .A1(d6_adj_5672[59]), 
          .B1(cout_adj_5179), .C1(n114_adj_5281), .D1(n14_adj_4680), .CIN(n15972), 
          .COUT(n15973), .S0(d7_71__N_1531_adj_5700[58]), .S1(d7_71__N_1531_adj_5700[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_23 (.A0(d6_adj_5672[56]), .B0(cout_adj_5179), 
          .C0(n123_adj_5284), .D0(n17_adj_4677), .A1(d6_adj_5672[57]), 
          .B1(cout_adj_5179), .C1(n120_adj_5283), .D1(n16_adj_4678), .CIN(n15971), 
          .COUT(n15972), .S0(d7_71__N_1531_adj_5700[56]), .S1(d7_71__N_1531_adj_5700[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_21 (.A0(d6_adj_5672[54]), .B0(cout_adj_5179), 
          .C0(n129_adj_5286), .D0(n19_adj_4675), .A1(d6_adj_5672[55]), 
          .B1(cout_adj_5179), .C1(n126_adj_5285), .D1(n18_adj_4676), .CIN(n15970), 
          .COUT(n15971), .S0(d7_71__N_1531_adj_5700[54]), .S1(d7_71__N_1531_adj_5700[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_19 (.A0(d6_adj_5672[52]), .B0(cout_adj_5179), 
          .C0(n135_adj_5288), .D0(n21_adj_4673), .A1(d6_adj_5672[53]), 
          .B1(cout_adj_5179), .C1(n132_adj_5287), .D1(n20_adj_4674), .CIN(n15969), 
          .COUT(n15970), .S0(d7_71__N_1531_adj_5700[52]), .S1(d7_71__N_1531_adj_5700[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_17 (.A0(d6_adj_5672[50]), .B0(cout_adj_5179), 
          .C0(n141_adj_5290), .D0(n23_adj_4671), .A1(d6_adj_5672[51]), 
          .B1(cout_adj_5179), .C1(n138_adj_5289), .D1(n22_adj_4672), .CIN(n15968), 
          .COUT(n15969), .S0(d7_71__N_1531_adj_5700[50]), .S1(d7_71__N_1531_adj_5700[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_37 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15846), .S0(n76));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1484_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_37.INJECT1_1 = "NO";
    LUT4 i3408_2_lut (.A(n250_adj_5638), .B(n17751), .Z(n2549)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3408_2_lut.init = 16'h8888;
    CCU2C _add_1_1637_add_4_6 (.A0(d_d7[39]), .B0(d7[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[40]), .B1(d7[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15922), .COUT(n15923), .S0(n174_adj_4921), .S1(n171_adj_4920));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_18 (.A0(d_d7[51]), .B0(d7[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[52]), .B1(d7[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15928), .COUT(n15929), .S0(n138_adj_4909), .S1(n135_adj_4908));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_18.INJECT1_1 = "NO";
    LUT4 i2264_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n253_adj_5639), .Z(n11953)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2264_3_lut_4_lut.init = 16'hf707;
    CCU2C _add_1_1472_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5216), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15574));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1472_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1472_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1472_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_4 (.A0(d_d7[37]), .B0(d7[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[38]), .B1(d7[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15921), .COUT(n15922), .S0(n180_adj_4923), .S1(n177_adj_4922));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1637_add_4_16 (.A0(d_d7[49]), .B0(d7[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[50]), .B1(d7[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15927), .COUT(n15928), .S0(n144_adj_4911), .S1(n141_adj_4910));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1637_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1637_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1637_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1637_add_4_16.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    CCU2C _add_1_1448_add_4_9 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n165_adj_5119), .D0(d1[42]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n162_adj_5118), .D1(d1[43]), .CIN(n15853), .COUT(n15854), 
          .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_9.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    CCU2C _add_1_1595_add_4_38 (.A0(d_d9_adj_5679[35]), .B0(d9_adj_5678[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15570), .S1(cout_adj_5089));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1595_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_38.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    CCU2C _add_1_1595_add_4_36 (.A0(d_d9_adj_5679[33]), .B0(d9_adj_5678[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[34]), .B1(d9_adj_5678[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15569), .COUT(n15570));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_36.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    CCU2C _add_1_1595_add_4_34 (.A0(d_d9_adj_5679[31]), .B0(d9_adj_5678[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[32]), .B1(d9_adj_5678[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15568), .COUT(n15569));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_32 (.A0(d_d9_adj_5679[29]), .B0(d9_adj_5678[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[30]), .B1(d9_adj_5678[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15567), .COUT(n15568));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_32.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i0 (.D(n321), .CK(clk_80mhz), .Q(phase_accum_adj_5658[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i0.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    CCU2C _add_1_1595_add_4_30 (.A0(d_d9_adj_5679[27]), .B0(d9_adj_5678[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[28]), .B1(d9_adj_5678[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15566), .COUT(n15567));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_28 (.A0(d_d9_adj_5679[25]), .B0(d9_adj_5678[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[26]), .B1(d9_adj_5678[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15565), .COUT(n15566));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_28.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    CCU2C _add_1_1466_add_4_19 (.A0(d7[52]), .B0(cout_adj_5088), .C0(n135_adj_4908), 
          .D0(n21_adj_4571), .A1(d7[53]), .B1(cout_adj_5088), .C1(n132_adj_4907), 
          .D1(n20_adj_4572), .CIN(n15910), .COUT(n15911), .S0(d8_71__N_1603[52]), 
          .S1(d8_71__N_1603[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_26 (.A0(d_d9_adj_5679[23]), .B0(d9_adj_5678[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[24]), .B1(d9_adj_5678[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15564), .COUT(n15565));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_26.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    CCU2C _add_1_1595_add_4_24 (.A0(d_d9_adj_5679[21]), .B0(d9_adj_5678[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[22]), .B1(d9_adj_5678[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15563), .COUT(n15564));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_22 (.A0(d_d9_adj_5679[19]), .B0(d9_adj_5678[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[20]), .B1(d9_adj_5678[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15562), .COUT(n15563));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_22.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i1 (.D(n126_adj_5178), .CK(CIC1_out_clkSin), .Q(ISquare[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i1.GSR = "ENABLED";
    CCU2C _add_1_1466_add_4_17 (.A0(d7[50]), .B0(cout_adj_5088), .C0(n141_adj_4910), 
          .D0(n23_adj_4836), .A1(d7[51]), .B1(cout_adj_5088), .C1(n138_adj_4909), 
          .D1(n22_adj_4570), .CIN(n15909), .COUT(n15910), .S0(d8_71__N_1603[50]), 
          .S1(d8_71__N_1603[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_20 (.A0(d_d9_adj_5679[17]), .B0(d9_adj_5678[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[18]), .B1(d9_adj_5678[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15561), .COUT(n15562));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_21 (.A0(d4_adj_5670[54]), .B0(cout_adj_5137), 
          .C0(n129), .D0(d5_adj_5671[54]), .A1(d4_adj_5670[55]), .B1(cout_adj_5137), 
          .C1(n126), .D1(d5_adj_5671[55]), .CIN(n15784), .COUT(n15785), 
          .S0(d5_71__N_706_adj_5687[54]), .S1(d5_71__N_706_adj_5687[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_19 (.A0(d4_adj_5670[52]), .B0(cout_adj_5137), 
          .C0(n135), .D0(d5_adj_5671[52]), .A1(d4_adj_5670[53]), .B1(cout_adj_5137), 
          .C1(n132), .D1(d5_adj_5671[53]), .CIN(n15783), .COUT(n15784), 
          .S0(d5_71__N_706_adj_5687[52]), .S1(d5_71__N_706_adj_5687[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_19.INJECT1_1 = "NO";
    LUT4 i2254_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n271_adj_5645), 
         .Z(n11943)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2254_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1595_add_4_18 (.A0(d_d9_adj_5679[15]), .B0(d9_adj_5678[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[16]), .B1(d9_adj_5678[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15560), .COUT(n15561));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_7 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n171_adj_5121), .D0(d1[40]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n168_adj_5120), .D1(d1[41]), .CIN(n15852), .COUT(n15853), 
          .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_15 (.A0(d7[48]), .B0(cout_adj_5088), .C0(n147_adj_4912), 
          .D0(n25), .A1(d7[49]), .B1(cout_adj_5088), .C1(n144_adj_4911), 
          .D1(n24_adj_4812), .CIN(n15908), .COUT(n15909), .S0(d8_71__N_1603[48]), 
          .S1(d8_71__N_1603[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_15.INJECT1_1 = "NO";
    LUT4 i2260_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n259_adj_5641), .Z(n11949)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2260_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_4_lut_then_4_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[2]), .C(MYLED_0_6), 
         .D(o_Rx_Byte[0]), .Z(n17647)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_4_lut_then_4_lut.init = 16'h4440;
    LUT4 i1_4_lut_else_4_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[2]), .C(MYLED_0_6), 
         .D(o_Rx_Byte[0]), .Z(n17646)) /* synthesis lut_function=(!(A+!(B (C)+!B !((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_4_lut_else_4_lut.init = 16'h4050;
    CCU2C _add_1_1439_add_4_28 (.A0(d4_adj_5670[26]), .B0(d3_adj_5669[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[27]), .B1(d3_adj_5669[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15993), .COUT(n15994), .S0(d4_71__N_634_adj_5686[26]), 
          .S1(d4_71__N_634_adj_5686[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_36 (.A0(d_d6_adj_5673[69]), .B0(d6_adj_5672[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[70]), .B1(d6_adj_5672[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16187), .COUT(n16188), .S0(n84_adj_5271), 
          .S1(n81_adj_5270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_36.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(o_Rx_Byte[4]), .B(n17632), .C(o_Rx_Byte[3]), 
         .D(o_Rx_Byte[2]), .Z(n16818)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_3_lut_rep_160 (.A(o_Rx_Byte[4]), .B(n17634), .C(o_Rx_Byte[0]), 
         .Z(n17629)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_3_lut_rep_160.init = 16'h8080;
    CCU2C _add_1_1439_add_4_26 (.A0(d4_adj_5670[24]), .B0(d3_adj_5669[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[25]), .B1(d3_adj_5669[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15992), .COUT(n15993), .S0(d4_71__N_634_adj_5686[24]), 
          .S1(d4_71__N_634_adj_5686[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_24 (.A0(d4_adj_5670[22]), .B0(d3_adj_5669[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[23]), .B1(d3_adj_5669[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15991), .COUT(n15992), .S0(d4_71__N_634_adj_5686[22]), 
          .S1(d4_71__N_634_adj_5686[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_24.INJECT1_1 = "NO";
    LUT4 i2804_2_lut_3_lut (.A(n12378), .B(n17633), .C(n17751), .Z(n12511)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i2804_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i5155_2_lut (.A(d2[0]), .B(d1[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5155_2_lut.init = 16'h6666;
    CCU2C _add_1_1490_add_4_17 (.A0(d4_adj_5670[50]), .B0(cout_adj_5137), 
          .C0(n141), .D0(d5_adj_5671[50]), .A1(d4_adj_5670[51]), .B1(cout_adj_5137), 
          .C1(n138), .D1(d5_adj_5671[51]), .CIN(n15782), .COUT(n15783), 
          .S0(d5_71__N_706_adj_5687[50]), .S1(d5_71__N_706_adj_5687[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_17.INJECT1_1 = "NO";
    LUT4 i5153_2_lut (.A(d3[0]), .B(d2[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5153_2_lut.init = 16'h6666;
    LUT4 i6166_4_lut_rep_208 (.A(n16740), .B(n17632), .C(n17648), .D(n17449), 
         .Z(n17784)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i6166_4_lut_rep_208.init = 16'h3032;
    CCU2C _add_1_1478_add_4_15 (.A0(d6_adj_5672[48]), .B0(cout_adj_5179), 
          .C0(n147_adj_5292), .D0(n25_adj_4669), .A1(d6_adj_5672[49]), 
          .B1(cout_adj_5179), .C1(n144_adj_5291), .D1(n24_adj_4670), .CIN(n15967), 
          .COUT(n15968), .S0(d7_71__N_1531_adj_5700[48]), .S1(d7_71__N_1531_adj_5700[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_15 (.A0(d4_adj_5670[48]), .B0(cout_adj_5137), 
          .C0(n147), .D0(d5_adj_5671[48]), .A1(d4_adj_5670[49]), .B1(cout_adj_5137), 
          .C1(n144), .D1(d5_adj_5671[49]), .CIN(n15781), .COUT(n15782), 
          .S0(d5_71__N_706_adj_5687[48]), .S1(d5_71__N_706_adj_5687[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_15.INJECT1_1 = "NO";
    LUT4 i6166_4_lut_rep_209 (.A(n16740), .B(n17632), .C(n17648), .D(n17449), 
         .Z(clk_80mhz_enable_1460)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i6166_4_lut_rep_209.init = 16'h3032;
    CCU2C _add_1_1595_add_4_16 (.A0(d_d9_adj_5679[13]), .B0(d9_adj_5678[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[14]), .B1(d9_adj_5678[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15559), .COUT(n15560));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_11 (.A0(d6_adj_5672[44]), .B0(cout_adj_5179), 
          .C0(n159_adj_5296), .D0(n29_adj_4665), .A1(d6_adj_5672[45]), 
          .B1(cout_adj_5179), .C1(n156_adj_5295), .D1(n28_adj_4666), .CIN(n15965), 
          .COUT(n15966), .S0(d7_71__N_1531_adj_5700[44]), .S1(d7_71__N_1531_adj_5700[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_9 (.A0(d6_adj_5672[42]), .B0(cout_adj_5179), 
          .C0(n165_adj_5298), .D0(n31_adj_4663), .A1(d6_adj_5672[43]), 
          .B1(cout_adj_5179), .C1(n162_adj_5297), .D1(n30_adj_4664), .CIN(n15964), 
          .COUT(n15965), .S0(d7_71__N_1531_adj_5700[42]), .S1(d7_71__N_1531_adj_5700[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_9.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i0 (.D(n323), .SP(clk_80mhz_enable_45), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1490_add_4_13 (.A0(d4_adj_5670[46]), .B0(cout_adj_5137), 
          .C0(n153), .D0(d5_adj_5671[46]), .A1(d4_adj_5670[47]), .B1(cout_adj_5137), 
          .C1(n150), .D1(d5_adj_5671[47]), .CIN(n15780), .COUT(n15781), 
          .S0(d5_71__N_706_adj_5687[46]), .S1(d5_71__N_706_adj_5687[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_13.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i0 (.D(o_Rx_Byte1[0]), .CK(clk_80mhz), .Q(o_Rx_Byte[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1S3AX _add_1_1649_i7 (.D(cout_adj_4998), .CK(clk_80mhz), .Q(PWMOutP4_c));
    defparam _add_1_1649_i7.GSR = "ENABLED";
    OB MYLED_pad_6 (.I(MYLED_0_6), .O(MYLED[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    CCU2C _add_1_1490_add_4_11 (.A0(d4_adj_5670[44]), .B0(cout_adj_5137), 
          .C0(n159), .D0(d5_adj_5671[44]), .A1(d4_adj_5670[45]), .B1(cout_adj_5137), 
          .C1(n156), .D1(d5_adj_5671[45]), .CIN(n15779), .COUT(n15780), 
          .S0(d5_71__N_706_adj_5687[44]), .S1(d5_71__N_706_adj_5687[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_9 (.A0(d4_adj_5670[42]), .B0(cout_adj_5137), 
          .C0(n165_adj_2768), .D0(d5_adj_5671[42]), .A1(d4_adj_5670[43]), 
          .B1(cout_adj_5137), .C1(n162), .D1(d5_adj_5671[43]), .CIN(n15778), 
          .COUT(n15779), .S0(d5_71__N_706_adj_5687[42]), .S1(d5_71__N_706_adj_5687[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_7 (.A0(d4_adj_5670[40]), .B0(cout_adj_5137), 
          .C0(n171_adj_2766), .D0(d5_adj_5671[40]), .A1(d4_adj_5670[41]), 
          .B1(cout_adj_5137), .C1(n168_adj_2767), .D1(d5_adj_5671[41]), 
          .CIN(n15777), .COUT(n15778), .S0(d5_71__N_706_adj_5687[40]), 
          .S1(d5_71__N_706_adj_5687[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_5 (.A0(d4_adj_5670[38]), .B0(cout_adj_5137), 
          .C0(n177_adj_2764), .D0(d5_adj_5671[38]), .A1(d4_adj_5670[39]), 
          .B1(cout_adj_5137), .C1(n174_adj_2765), .D1(d5_adj_5671[39]), 
          .CIN(n15776), .COUT(n15777), .S0(d5_71__N_706_adj_5687[38]), 
          .S1(d5_71__N_706_adj_5687[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_3 (.A0(d4_adj_5670[36]), .B0(cout_adj_5137), 
          .C0(n183), .D0(d5_adj_5671[36]), .A1(d4_adj_5670[37]), .B1(cout_adj_5137), 
          .C1(n180_adj_2763), .D1(d5_adj_5671[37]), .CIN(n15775), .COUT(n15776), 
          .S0(d5_71__N_706_adj_5687[36]), .S1(d5_71__N_706_adj_5687[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_13 (.A0(d6_adj_5672[46]), .B0(cout_adj_5179), 
          .C0(n153_adj_5294), .D0(n27_adj_4667), .A1(d6_adj_5672[47]), 
          .B1(cout_adj_5179), .C1(n150_adj_5293), .D1(n26_adj_4668), .CIN(n15966), 
          .COUT(n15967), .S0(d7_71__N_1531_adj_5700[46]), .S1(d7_71__N_1531_adj_5700[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5137), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15775));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1490_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1490_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_34 (.A0(d_d6_adj_5673[67]), .B0(d6_adj_5672[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[68]), .B1(d6_adj_5672[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16186), .COUT(n16187), .S0(n90_adj_5273), 
          .S1(n87_adj_5272));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_34.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_159_3_lut (.A(o_Rx_Byte[6]), .B(n17638), .C(o_Rx_Byte[4]), 
         .Z(n17628)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_2_lut_rep_159_3_lut.init = 16'hfdfd;
    CCU2C _add_1_1574_add_4_38 (.A0(d4_adj_5670[71]), .B0(d3_adj_5669[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15771), .S0(n78_adj_4565));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1574_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_36 (.A0(d4_adj_5670[69]), .B0(d3_adj_5669[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[70]), .B1(d3_adj_5669[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15770), .COUT(n15771), .S0(n84_adj_4563), 
          .S1(n81_adj_4564));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_14 (.A0(d5_adj_5671[12]), .B0(d4_adj_5670[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[13]), .B1(d4_adj_5670[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15945), .COUT(n15946), .S0(d5_71__N_706_adj_5687[12]), 
          .S1(d5_71__N_706_adj_5687[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_34 (.A0(d4_adj_5670[67]), .B0(d3_adj_5669[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[68]), .B1(d3_adj_5669[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15769), .COUT(n15770), .S0(n90_adj_4561), 
          .S1(n87_adj_4562));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_32 (.A0(d_d6_adj_5673[65]), .B0(d6_adj_5672[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[66]), .B1(d6_adj_5672[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16185), .COUT(n16186), .S0(n96_adj_5275), 
          .S1(n93_adj_5274));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_32 (.A0(d4_adj_5670[65]), .B0(d3_adj_5669[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[66]), .B1(d3_adj_5669[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15768), .COUT(n15769), .S0(n96_adj_4559), 
          .S1(n93_adj_4560));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_30 (.A0(d4_adj_5670[63]), .B0(d3_adj_5669[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[64]), .B1(d3_adj_5669[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15767), .COUT(n15768), .S0(n102_adj_4557), 
          .S1(n99_adj_4558));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_22 (.A0(d4_adj_5670[20]), .B0(d3_adj_5669[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[21]), .B1(d3_adj_5669[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15990), .COUT(n15991), .S0(d4_71__N_634_adj_5686[20]), 
          .S1(d4_71__N_634_adj_5686[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_28 (.A0(d4_adj_5670[61]), .B0(d3_adj_5669[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[62]), .B1(d3_adj_5669[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15766), .COUT(n15767), .S0(n108_adj_4555), 
          .S1(n105_adj_4556));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_26 (.A0(d4_adj_5670[59]), .B0(d3_adj_5669[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[60]), .B1(d3_adj_5669[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15765), .COUT(n15766), .S0(n114_adj_4553), 
          .S1(n111_adj_4554));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_24 (.A0(d4_adj_5670[57]), .B0(d3_adj_5669[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[58]), .B1(d3_adj_5669[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15764), .COUT(n15765), .S0(n120_adj_4551), 
          .S1(n117_adj_4552));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_24.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_165 (.A(n12378), .B(n17750), .C(MYLED_0_6), .Z(n17634)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_3_lut_rep_165.init = 16'h0202;
    CCU2C _add_1_1574_add_4_22 (.A0(d4_adj_5670[55]), .B0(d3_adj_5669[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[56]), .B1(d3_adj_5669[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15763), .COUT(n15764), .S0(n126_adj_4549), 
          .S1(n123_adj_4550));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_20 (.A0(d4_adj_5670[53]), .B0(d3_adj_5669[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[54]), .B1(d3_adj_5669[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15762), .COUT(n15763), .S0(n132_adj_4547), 
          .S1(n129_adj_4548));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_20 (.A0(d4_adj_5670[18]), .B0(d3_adj_5669[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[19]), .B1(d3_adj_5669[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15989), .COUT(n15990), .S0(d4_71__N_634_adj_5686[18]), 
          .S1(d4_71__N_634_adj_5686[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1439_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_18 (.A0(d4_adj_5670[51]), .B0(d3_adj_5669[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[52]), .B1(d3_adj_5669[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15761), .COUT(n15762), .S0(n138_adj_4545), 
          .S1(n135_adj_4546));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_16 (.A0(d4_adj_5670[49]), .B0(d3_adj_5669[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[50]), .B1(d3_adj_5669[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15760), .COUT(n15761), .S0(n144_adj_4543), 
          .S1(n141_adj_4544));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_14 (.A0(d4_adj_5670[47]), .B0(d3_adj_5669[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[48]), .B1(d3_adj_5669[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15759), .COUT(n15760), .S0(n150_adj_4541), 
          .S1(n147_adj_4542));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_14.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_162_4_lut (.A(n12378), .B(n17750), .C(MYLED_0_6), 
         .D(n17637), .Z(n17631)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_2_lut_rep_162_4_lut.init = 16'h0200;
    CCU2C _add_1_1574_add_4_12 (.A0(d4_adj_5670[45]), .B0(d3_adj_5669[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[46]), .B1(d3_adj_5669[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15758), .COUT(n15759), .S0(n156_adj_4520), 
          .S1(n153_adj_4540));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_30 (.A0(d_d6_adj_5673[63]), .B0(d6_adj_5672[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[64]), .B1(d6_adj_5672[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16184), .COUT(n16185), .S0(n102_adj_5277), 
          .S1(n99_adj_5276));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_10 (.A0(d4_adj_5670[43]), .B0(d3_adj_5669[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[44]), .B1(d3_adj_5669[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15757), .COUT(n15758), .S0(n162_adj_3854), 
          .S1(n159_adj_3855));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_36 (.A0(d5_adj_5671[34]), .B0(d4_adj_5670[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[35]), .B1(d4_adj_5670[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15956), .COUT(n15957), .S0(d5_71__N_706_adj_5687[34]), 
          .S1(d5_71__N_706_adj_5687[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_18 (.A0(d5_adj_5671[16]), .B0(d4_adj_5670[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[17]), .B1(d4_adj_5670[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15947), .COUT(n15948), .S0(d5_71__N_706_adj_5687[16]), 
          .S1(d5_71__N_706_adj_5687[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_30 (.A0(d5_adj_5671[28]), .B0(d4_adj_5670[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[29]), .B1(d4_adj_5670[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15953), .COUT(n15954), .S0(d5_71__N_706_adj_5687[28]), 
          .S1(d5_71__N_706_adj_5687[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1442_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1442_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1442_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_8 (.A0(d4_adj_5670[41]), .B0(d3_adj_5669[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[42]), .B1(d3_adj_5669[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15756), .COUT(n15757), .S0(n168), 
          .S1(n165));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1574_add_4_6 (.A0(d4_adj_5670[39]), .B0(d3_adj_5669[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[40]), .B1(d3_adj_5669[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15755), .COUT(n15756), .S0(n174), 
          .S1(n171));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_6.INJECT1_1 = "NO";
    OB MYLED_pad_7 (.I(GND_net), .O(MYLED[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    CCU2C _add_1_1625_add_4_28 (.A0(d_d6_adj_5673[61]), .B0(d6_adj_5672[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[62]), .B1(d6_adj_5672[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16183), .COUT(n16184), .S0(n108_adj_5279), 
          .S1(n105_adj_5278));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_28.INJECT1_1 = "NO";
    OB o_Tx_Serial_pad (.I(GND_net), .O(o_Tx_Serial));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(49[11:22])
    \uart_rx(CLKS_PER_BIT=87)  uart_rx1 (.clk_80mhz(clk_80mhz), .i_Rx_Serial_c(i_Rx_Serial_c), 
            .o_Rx_Byte1({o_Rx_Byte1}), .o_Rx_DV1(o_Rx_DV1), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(229[32] 234[2])
    CCU2C _add_1_1574_add_4_4 (.A0(d4_adj_5670[37]), .B0(d3_adj_5669[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5670[38]), .B1(d3_adj_5669[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15754), .COUT(n15755), .S0(n180), 
          .S1(n177));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1574_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_4.INJECT1_1 = "NO";
    OB MYLED_pad_5 (.I(MYLED_0_5), .O(MYLED[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    LUT4 i5158_2_lut (.A(d4[0]), .B(d3[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5158_2_lut.init = 16'h6666;
    FD1S3AX o_Rx_Byte_i7 (.D(o_Rx_Byte1[7]), .CK(clk_80mhz), .Q(o_Rx_Byte[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i6 (.D(o_Rx_Byte1[6]), .CK(clk_80mhz), .Q(o_Rx_Byte[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i5 (.D(o_Rx_Byte1[5]), .CK(clk_80mhz), .Q(o_Rx_Byte[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i4 (.D(o_Rx_Byte1[4]), .CK(clk_80mhz), .Q(o_Rx_Byte[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i3 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(o_Rx_Byte[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i2 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(o_Rx_Byte[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i1 (.D(o_Rx_Byte1[1]), .CK(clk_80mhz), .Q(MYLED_0_6));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    CCU2C _add_1_1574_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4_adj_5670[36]), .B1(d3_adj_5669[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15754), .S1(n183_adj_4539));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1574_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1574_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1574_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1574_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_38 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15753), .S0(n78_adj_5037));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1583_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_38.INJECT1_1 = "NO";
    LUT4 n2660_bdd_4_lut_6220 (.A(o_Rx_Byte[0]), .B(o_Rx_Byte[4]), .C(MYLED_0_6), 
         .D(o_Rx_Byte[2]), .Z(n17572)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B+!(C)))) */ ;
    defparam n2660_bdd_4_lut_6220.init = 16'h301a;
    CCU2C ISquare_add_4_10 (.A0(MultResult2[8]), .B0(MultResult1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[9]), .B1(MultResult1[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15798), .COUT(n15799), .S0(n102_adj_5170), 
          .S1(n99_adj_5169));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_10.INIT0 = 16'h666a;
    defparam ISquare_add_4_10.INIT1 = 16'h666a;
    defparam ISquare_add_4_10.INJECT1_0 = "NO";
    defparam ISquare_add_4_10.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_8 (.A0(MultResult2[6]), .B0(MultResult1[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[7]), .B1(MultResult1[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15797), .COUT(n15798), .S0(n108_adj_5172), 
          .S1(n105_adj_5171));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_8.INIT0 = 16'h666a;
    defparam ISquare_add_4_8.INIT1 = 16'h666a;
    defparam ISquare_add_4_8.INJECT1_0 = "NO";
    defparam ISquare_add_4_8.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_168 (.A(o_Rx_Byte[0]), .B(o_Rx_Byte[4]), .Z(n17637)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_2_lut_rep_168.init = 16'h2222;
    OB MYLED_pad_4 (.I(MYLED_0_4), .O(MYLED[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    OB MYLED_pad_3 (.I(MYLED_0_3), .O(MYLED[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    OB MYLED_pad_2 (.I(MYLED_0_2), .O(MYLED[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    OB MYLED_pad_1 (.I(MYLED_0_1), .O(MYLED[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    OB MYLED_pad_0 (.I(MYLED_0_0), .O(MYLED[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(50[18:23])
    OB XOut_pad (.I(GND_net), .O(XOut));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(54[9:13])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(56[9:16])
    OB PWMOut_pad (.I(PWMOutP4_c), .O(PWMOut));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(57[9:15])
    OB PWMOutP1_pad (.I(PWMOutP4_c), .O(PWMOutP1));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(58[9:17])
    OB PWMOutP2_pad (.I(PWMOutP4_c), .O(PWMOutP2));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(59[9:17])
    OB PWMOutP3_pad (.I(PWMOutP4_c), .O(PWMOutP3));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(60[9:17])
    OB PWMOutP4_pad (.I(PWMOutP4_c), .O(PWMOutP4));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(61[9:17])
    OB PWMOutN1_pad (.I(PWMOutN4_c), .O(PWMOutN1));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(62[9:17])
    OB PWMOutN2_pad (.I(PWMOutN4_c), .O(PWMOutN2));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(63[9:17])
    OB PWMOutN3_pad (.I(PWMOutN4_c), .O(PWMOutN3));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(64[9:17])
    OB PWMOutN4_pad (.I(PWMOutN4_c), .O(PWMOutN4));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(65[9:17])
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(66[9:15])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(67[9:16])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(68[9:23])
    IB osc_clk_pad (.I(osc_clk), .O(osc_clk_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(47[13:20])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(48[13:24])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(55[9:13])
    CCU2C _add_1_1466_add_4_13 (.A0(d7[46]), .B0(cout_adj_5088), .C0(n153_adj_4914), 
          .D0(n27), .A1(d7[47]), .B1(cout_adj_5088), .C1(n150_adj_4913), 
          .D1(n26), .CIN(n15907), .COUT(n15908), .S0(d8_71__N_1603[46]), 
          .S1(d8_71__N_1603[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_11 (.A0(d7[44]), .B0(cout_adj_5088), .C0(n159_adj_4916), 
          .D0(n29), .A1(d7[45]), .B1(cout_adj_5088), .C1(n156_adj_4915), 
          .D1(n28), .CIN(n15906), .COUT(n15907), .S0(d8_71__N_1603[44]), 
          .S1(d8_71__N_1603[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_9 (.A0(d7[42]), .B0(cout_adj_5088), .C0(n165_adj_4918), 
          .D0(n31), .A1(d7[43]), .B1(cout_adj_5088), .C1(n162_adj_4917), 
          .D1(n30), .CIN(n15905), .COUT(n15906), .S0(d8_71__N_1603[42]), 
          .S1(d8_71__N_1603[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_7 (.A0(d7[40]), .B0(cout_adj_5088), .C0(n171_adj_4920), 
          .D0(n33_adj_4697), .A1(d7[41]), .B1(cout_adj_5088), .C1(n168_adj_4919), 
          .D1(n32), .CIN(n15904), .COUT(n15905), .S0(d8_71__N_1603[40]), 
          .S1(d8_71__N_1603[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(o_Rx_Byte[0]), .B(o_Rx_Byte[4]), .C(MYLED_0_6), 
         .D(n17751), .Z(n16930)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_3_lut_4_lut.init = 16'h2000;
    CCU2C _add_1_1466_add_4_5 (.A0(d7[38]), .B0(cout_adj_5088), .C0(n177_adj_4922), 
          .D0(n35_adj_4695), .A1(d7[39]), .B1(cout_adj_5088), .C1(n174_adj_4921), 
          .D1(n34_adj_4696), .CIN(n15903), .COUT(n15904), .S0(d8_71__N_1603[38]), 
          .S1(d8_71__N_1603[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_3 (.A0(d7[36]), .B0(cout_adj_5088), .C0(n183_adj_4924), 
          .D0(n37_adj_4688), .A1(d7[37]), .B1(cout_adj_5088), .C1(n180_adj_4923), 
          .D1(n36_adj_4694), .CIN(n15902), .COUT(n15903), .S0(d8_71__N_1603[36]), 
          .S1(d8_71__N_1603[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1466_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1466_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5088), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15902));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1466_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1466_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1466_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_1.INJECT1_1 = "NO";
    LUT4 i5157_2_lut (.A(d5[0]), .B(d4[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5157_2_lut.init = 16'h6666;
    CCU2C _add_1_1445_add_4_17 (.A0(count_adj_5682[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15898), .S0(n36_adj_5138));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1445_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_15 (.A0(count_adj_5682[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15897), .COUT(n15898), .S0(n42_adj_5140), 
          .S1(n39_adj_5139));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_13 (.A0(count_adj_5682[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15896), .COUT(n15897), .S0(n48_adj_5142), 
          .S1(n45_adj_5141));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_11 (.A0(count_adj_5682[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15895), .COUT(n15896), .S0(n54_adj_5144), 
          .S1(n51_adj_5143));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_9 (.A0(count_adj_5682[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15894), .COUT(n15895), .S0(n60_adj_5146), 
          .S1(n57_adj_5145));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_7 (.A0(count_adj_5682[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15893), .COUT(n15894), .S0(n66_adj_5148), 
          .S1(n63_adj_5147));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_5 (.A0(count_adj_5682[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15892), .COUT(n15893), .S0(n72_adj_5150), 
          .S1(n69_adj_5149));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_3 (.A0(count_adj_5682[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5682[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15891), .COUT(n15892), .S0(n78_adj_5152), 
          .S1(n75_adj_5151));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1445_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1445_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_adj_5682[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15891), .S1(n81_adj_5153));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1445_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1445_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1445_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_37 (.A0(d_tmp_adj_5665[70]), .B0(cout_adj_5420), 
          .C0(n81_adj_5053), .D0(n3_adj_2761), .A1(d_tmp_adj_5665[71]), 
          .B1(cout_adj_5420), .C1(n78_adj_5052), .D1(n2_adj_2762), .CIN(n15889), 
          .S0(d6_71__N_1459_adj_5699[70]), .S1(d6_71__N_1459_adj_5699[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_35 (.A0(d_tmp_adj_5665[68]), .B0(cout_adj_5420), 
          .C0(n87_adj_5055), .D0(n5_adj_2759), .A1(d_tmp_adj_5665[69]), 
          .B1(cout_adj_5420), .C1(n84_adj_5054), .D1(n4_adj_2760), .CIN(n15888), 
          .COUT(n15889), .S0(d6_71__N_1459_adj_5699[68]), .S1(d6_71__N_1459_adj_5699[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_33 (.A0(d_tmp_adj_5665[66]), .B0(cout_adj_5420), 
          .C0(n93_adj_5057), .D0(n7_adj_2757), .A1(d_tmp_adj_5665[67]), 
          .B1(cout_adj_5420), .C1(n90_adj_5056), .D1(n6_adj_2758), .CIN(n15887), 
          .COUT(n15888), .S0(d6_71__N_1459_adj_5699[66]), .S1(d6_71__N_1459_adj_5699[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_31 (.A0(d_tmp_adj_5665[64]), .B0(cout_adj_5420), 
          .C0(n99_adj_5059), .D0(n9), .A1(d_tmp_adj_5665[65]), .B1(cout_adj_5420), 
          .C1(n96_adj_5058), .D1(n8), .CIN(n15886), .COUT(n15887), .S0(d6_71__N_1459_adj_5699[64]), 
          .S1(d6_71__N_1459_adj_5699[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_29 (.A0(d_tmp_adj_5665[62]), .B0(cout_adj_5420), 
          .C0(n105_adj_5061), .D0(n11), .A1(d_tmp_adj_5665[63]), .B1(cout_adj_5420), 
          .C1(n102_adj_5060), .D1(n10), .CIN(n15885), .COUT(n15886), 
          .S0(d6_71__N_1459_adj_5699[62]), .S1(d6_71__N_1459_adj_5699[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_27 (.A0(d_tmp_adj_5665[60]), .B0(cout_adj_5420), 
          .C0(n111_adj_5063), .D0(n13), .A1(d_tmp_adj_5665[61]), .B1(cout_adj_5420), 
          .C1(n108_adj_5062), .D1(n12), .CIN(n15884), .COUT(n15885), 
          .S0(d6_71__N_1459_adj_5699[60]), .S1(d6_71__N_1459_adj_5699[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_25 (.A0(d_tmp_adj_5665[58]), .B0(cout_adj_5420), 
          .C0(n117_adj_5065), .D0(n15), .A1(d_tmp_adj_5665[59]), .B1(cout_adj_5420), 
          .C1(n114_adj_5064), .D1(n14), .CIN(n15883), .COUT(n15884), 
          .S0(d6_71__N_1459_adj_5699[58]), .S1(d6_71__N_1459_adj_5699[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_25.INJECT1_1 = "NO";
    LUT4 i2244_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n289_adj_5651), .Z(n11933)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2244_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1481_add_4_23 (.A0(d_tmp_adj_5665[56]), .B0(cout_adj_5420), 
          .C0(n123_adj_5067), .D0(n17), .A1(d_tmp_adj_5665[57]), .B1(cout_adj_5420), 
          .C1(n120_adj_5066), .D1(n16), .CIN(n15882), .COUT(n15883), 
          .S0(d6_71__N_1459_adj_5699[56]), .S1(d6_71__N_1459_adj_5699[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_21 (.A0(d_tmp_adj_5665[54]), .B0(cout_adj_5420), 
          .C0(n129_adj_5069), .D0(n19), .A1(d_tmp_adj_5665[55]), .B1(cout_adj_5420), 
          .C1(n126_adj_5068), .D1(n18), .CIN(n15881), .COUT(n15882), 
          .S0(d6_71__N_1459_adj_5699[54]), .S1(d6_71__N_1459_adj_5699[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_19 (.A0(d_tmp_adj_5665[52]), .B0(cout_adj_5420), 
          .C0(n135_adj_5071), .D0(n21), .A1(d_tmp_adj_5665[53]), .B1(cout_adj_5420), 
          .C1(n132_adj_5070), .D1(n20), .CIN(n15880), .COUT(n15881), 
          .S0(d6_71__N_1459_adj_5699[52]), .S1(d6_71__N_1459_adj_5699[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_17 (.A0(d_tmp_adj_5665[50]), .B0(cout_adj_5420), 
          .C0(n141_adj_5073), .D0(n23), .A1(d_tmp_adj_5665[51]), .B1(cout_adj_5420), 
          .C1(n138_adj_5072), .D1(n22), .CIN(n15879), .COUT(n15880), 
          .S0(d6_71__N_1459_adj_5699[50]), .S1(d6_71__N_1459_adj_5699[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_15 (.A0(d_tmp_adj_5665[48]), .B0(cout_adj_5420), 
          .C0(n147_adj_5075), .D0(n25_adj_2756), .A1(d_tmp_adj_5665[49]), 
          .B1(cout_adj_5420), .C1(n144_adj_5074), .D1(n24), .CIN(n15878), 
          .COUT(n15879), .S0(d6_71__N_1459_adj_5699[48]), .S1(d6_71__N_1459_adj_5699[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_13 (.A0(d_tmp_adj_5665[46]), .B0(cout_adj_5420), 
          .C0(n153_adj_5077), .D0(n27_adj_2754), .A1(d_tmp_adj_5665[47]), 
          .B1(cout_adj_5420), .C1(n150_adj_5076), .D1(n26_adj_2755), .CIN(n15877), 
          .COUT(n15878), .S0(d6_71__N_1459_adj_5699[46]), .S1(d6_71__N_1459_adj_5699[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_11 (.A0(d_tmp_adj_5665[44]), .B0(cout_adj_5420), 
          .C0(n159_adj_5079), .D0(n29_adj_2752), .A1(d_tmp_adj_5665[45]), 
          .B1(cout_adj_5420), .C1(n156_adj_5078), .D1(n28_adj_2753), .CIN(n15876), 
          .COUT(n15877), .S0(d6_71__N_1459_adj_5699[44]), .S1(d6_71__N_1459_adj_5699[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_9 (.A0(d_tmp_adj_5665[42]), .B0(cout_adj_5420), 
          .C0(n165_adj_5081), .D0(n31_adj_2750), .A1(d_tmp_adj_5665[43]), 
          .B1(cout_adj_5420), .C1(n162_adj_5080), .D1(n30_adj_2751), .CIN(n15875), 
          .COUT(n15876), .S0(d6_71__N_1459_adj_5699[42]), .S1(d6_71__N_1459_adj_5699[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_7 (.A0(d_tmp_adj_5665[40]), .B0(cout_adj_5420), 
          .C0(n171_adj_5083), .D0(n33), .A1(d_tmp_adj_5665[41]), .B1(cout_adj_5420), 
          .C1(n168_adj_5082), .D1(n32_adj_2749), .CIN(n15874), .COUT(n15875), 
          .S0(d6_71__N_1459_adj_5699[40]), .S1(d6_71__N_1459_adj_5699[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_5 (.A0(d_tmp_adj_5665[38]), .B0(cout_adj_5420), 
          .C0(n177_adj_5085), .D0(n35), .A1(d_tmp_adj_5665[39]), .B1(cout_adj_5420), 
          .C1(n174_adj_5084), .D1(n34), .CIN(n15873), .COUT(n15874), 
          .S0(d6_71__N_1459_adj_5699[38]), .S1(d6_71__N_1459_adj_5699[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_3 (.A0(d_tmp_adj_5665[36]), .B0(cout_adj_5420), 
          .C0(n183_adj_5087), .D0(n37), .A1(d_tmp_adj_5665[37]), .B1(cout_adj_5420), 
          .C1(n180_adj_5086), .D1(n36), .CIN(n15872), .COUT(n15873), 
          .S0(d6_71__N_1459_adj_5699[36]), .S1(d6_71__N_1459_adj_5699[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1481_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1481_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5420), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15872));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1481_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1481_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1481_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_37 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n81_adj_5091), .D0(d1[70]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n78_adj_5090), .D1(d1[71]), .CIN(n15867), .S0(d1_71__N_418[70]), 
          .S1(d1_71__N_418[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_35 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n87_adj_5093), .D0(d1[68]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n84_adj_5092), .D1(d1[69]), .CIN(n15866), .COUT(n15867), 
          .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_33 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n93_adj_5095), .D0(d1[66]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n90_adj_5094), .D1(d1[67]), .CIN(n15865), .COUT(n15866), 
          .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_31 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n99_adj_5097), .D0(d1[64]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n96_adj_5096), .D1(d1[65]), .CIN(n15864), .COUT(n15865), 
          .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_29 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n105_adj_5099), .D0(d1[62]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n102_adj_5098), .D1(d1[63]), .CIN(n15863), .COUT(n15864), 
          .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_27 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n111_adj_5101), .D0(d1[60]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n108_adj_5100), .D1(d1[61]), .CIN(n15862), .COUT(n15863), 
          .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_27.INJECT1_1 = "NO";
    LUT4 i6127_3_lut (.A(o_Rx_Byte[3]), .B(n17784), .C(n13169), .Z(clk_80mhz_enable_1471)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;
    defparam i6127_3_lut.init = 16'hc4c4;
    CCU2C _add_1_1625_add_4_26 (.A0(d_d6_adj_5673[59]), .B0(d6_adj_5672[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[60]), .B1(d6_adj_5672[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16182), .COUT(n16183), .S0(n114_adj_5281), 
          .S1(n111_adj_5280));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_24 (.A0(d_d6_adj_5673[57]), .B0(d6_adj_5672[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[58]), .B1(d6_adj_5672[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16181), .COUT(n16182), .S0(n120_adj_5283), 
          .S1(n117_adj_5282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_22 (.A0(d_d6_adj_5673[55]), .B0(d6_adj_5672[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[56]), .B1(d6_adj_5672[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16180), .COUT(n16181), .S0(n126_adj_5285), 
          .S1(n123_adj_5284));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_20 (.A0(d_d6_adj_5673[53]), .B0(d6_adj_5672[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[54]), .B1(d6_adj_5672[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16179), .COUT(n16180), .S0(n132_adj_5287), 
          .S1(n129_adj_5286));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_18 (.A0(d_d6_adj_5673[51]), .B0(d6_adj_5672[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[52]), .B1(d6_adj_5672[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16178), .COUT(n16179), .S0(n138_adj_5289), 
          .S1(n135_adj_5288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_16 (.A0(d_d6_adj_5673[49]), .B0(d6_adj_5672[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[50]), .B1(d6_adj_5672[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16177), .COUT(n16178), .S0(n144_adj_5291), 
          .S1(n141_adj_5290));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_14 (.A0(d_d6_adj_5673[47]), .B0(d6_adj_5672[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[48]), .B1(d6_adj_5672[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16176), .COUT(n16177), .S0(n150_adj_5293), 
          .S1(n147_adj_5292));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_12 (.A0(d_d6_adj_5673[45]), .B0(d6_adj_5672[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[46]), .B1(d6_adj_5672[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16175), .COUT(n16176), .S0(n156_adj_5295), 
          .S1(n153_adj_5294));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_10 (.A0(d_d6_adj_5673[43]), .B0(d6_adj_5672[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[44]), .B1(d6_adj_5672[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16174), .COUT(n16175), .S0(n162_adj_5297), 
          .S1(n159_adj_5296));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_8 (.A0(d_d6_adj_5673[41]), .B0(d6_adj_5672[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[42]), .B1(d6_adj_5672[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16173), .COUT(n16174), .S0(n168_adj_5299), 
          .S1(n165_adj_5298));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_6 (.A0(d_d6_adj_5673[39]), .B0(d6_adj_5672[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[40]), .B1(d6_adj_5672[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16172), .COUT(n16173), .S0(n174_adj_5301), 
          .S1(n171_adj_5300));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_4 (.A0(d_d6_adj_5673[37]), .B0(d6_adj_5672[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[38]), .B1(d6_adj_5672[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16171), .COUT(n16172), .S0(n180_adj_5303), 
          .S1(n177_adj_5302));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1625_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1625_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5673[36]), .B1(d6_adj_5672[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16171), .S1(n183_adj_5304));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1625_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1625_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1625_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1625_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_38 (.A0(d_d8_adj_5677[71]), .B0(d8_adj_5676[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16170), .S0(n78));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1631_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_36 (.A0(d_d8_adj_5677[69]), .B0(d8_adj_5676[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[70]), .B1(d8_adj_5676[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16169), .COUT(n16170), .S0(n84), 
          .S1(n81));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_34 (.A0(d_d8_adj_5677[67]), .B0(d8_adj_5676[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[68]), .B1(d8_adj_5676[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16168), .COUT(n16169), .S0(n90), 
          .S1(n87));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_32 (.A0(d_d8_adj_5677[65]), .B0(d8_adj_5676[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[66]), .B1(d8_adj_5676[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16167), .COUT(n16168), .S0(n96_adj_4790), 
          .S1(n93_adj_4813));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_30 (.A0(d_d8_adj_5677[63]), .B0(d8_adj_5676[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[64]), .B1(d8_adj_5676[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16166), .COUT(n16167), .S0(n102_adj_4788), 
          .S1(n99_adj_4789));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_28 (.A0(d_d8_adj_5677[61]), .B0(d8_adj_5676[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[62]), .B1(d8_adj_5676[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16165), .COUT(n16166), .S0(n108_adj_4786), 
          .S1(n105_adj_4787));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_26 (.A0(d_d8_adj_5677[59]), .B0(d8_adj_5676[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[60]), .B1(d8_adj_5676[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16164), .COUT(n16165), .S0(n114_adj_4784), 
          .S1(n111_adj_4785));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_24 (.A0(d_d8_adj_5677[57]), .B0(d8_adj_5676[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[58]), .B1(d8_adj_5676[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16163), .COUT(n16164), .S0(n120_adj_4782), 
          .S1(n117_adj_4783));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_22 (.A0(d_d8_adj_5677[55]), .B0(d8_adj_5676[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[56]), .B1(d8_adj_5676[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16162), .COUT(n16163), .S0(n126_adj_4766), 
          .S1(n123_adj_4767));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_20 (.A0(d_d8_adj_5677[53]), .B0(d8_adj_5676[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[54]), .B1(d8_adj_5676[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16161), .COUT(n16162), .S0(n132_adj_4750), 
          .S1(n129_adj_4765));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_18 (.A0(d_d8_adj_5677[51]), .B0(d8_adj_5676[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[52]), .B1(d8_adj_5676[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16160), .COUT(n16161), .S0(n138_adj_4748), 
          .S1(n135_adj_4749));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_18.INJECT1_1 = "NO";
    LUT4 i2412_3_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(n17631), .C(n17633), 
         .D(n12378), .Z(n12108)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i2412_3_lut_4_lut_4_lut.init = 16'h5444;
    CCU2C _add_1_1631_add_4_16 (.A0(d_d8_adj_5677[49]), .B0(d8_adj_5676[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[50]), .B1(d8_adj_5676[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16159), .COUT(n16160), .S0(n144_adj_4746), 
          .S1(n141_adj_4747));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_14 (.A0(d_d8_adj_5677[47]), .B0(d8_adj_5676[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[48]), .B1(d8_adj_5676[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16158), .COUT(n16159), .S0(n150_adj_4744), 
          .S1(n147_adj_4745));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_12 (.A0(d_d8_adj_5677[45]), .B0(d8_adj_5676[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[46]), .B1(d8_adj_5676[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16157), .COUT(n16158), .S0(n156_adj_4742), 
          .S1(n153_adj_4743));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_10 (.A0(d_d8_adj_5677[43]), .B0(d8_adj_5676[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[44]), .B1(d8_adj_5676[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16156), .COUT(n16157), .S0(n162_adj_4740), 
          .S1(n159_adj_4741));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_10.INJECT1_1 = "NO";
    FD1P3AX CICGain__i2 (.D(MYLED_0_6), .SP(clk_80mhz_enable_1408), .CK(clk_80mhz), 
            .Q(CICGain[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam CICGain__i2.GSR = "ENABLED";
    CCU2C _add_1_1631_add_4_8 (.A0(d_d8_adj_5677[41]), .B0(d8_adj_5676[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[42]), .B1(d8_adj_5676[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16155), .COUT(n16156), .S0(n168_adj_4738), 
          .S1(n165_adj_4739));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_6 (.A0(d_d8_adj_5677[39]), .B0(d8_adj_5676[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[40]), .B1(d8_adj_5676[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16154), .COUT(n16155), .S0(n174_adj_4736), 
          .S1(n171_adj_4737));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_4 (.A0(d_d8_adj_5677[37]), .B0(d8_adj_5676[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[38]), .B1(d8_adj_5676[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16153), .COUT(n16154), .S0(n180_adj_4734), 
          .S1(n177_adj_4735));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1631_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_36 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15752), .COUT(n15753), .S0(n84_adj_5039), .S1(n81_adj_5038));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1631_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5677[36]), .B1(d8_adj_5676[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16153), .S1(n183_adj_4733));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1631_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1631_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1631_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1631_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_38 (.A0(d_d7_adj_5675[71]), .B0(d7_adj_5674[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16152), .S0(n78_adj_5305));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1628_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_38.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_20 (.A0(MultResult2[18]), .B0(MultResult1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[19]), .B1(MultResult1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15803), .COUT(n15804), .S0(n72_adj_5160), 
          .S1(n69_adj_5159));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_20.INIT0 = 16'h666a;
    defparam ISquare_add_4_20.INIT1 = 16'h666a;
    defparam ISquare_add_4_20.INJECT1_0 = "NO";
    defparam ISquare_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_34 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15751), .COUT(n15752), .S0(n90_adj_5041), .S1(n87_adj_5040));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_5 (.A0(d6_adj_5672[38]), .B0(cout_adj_5179), 
          .C0(n177_adj_5302), .D0(n35_adj_4659), .A1(d6_adj_5672[39]), 
          .B1(cout_adj_5179), .C1(n174_adj_5301), .D1(n34_adj_4660), .CIN(n15962), 
          .COUT(n15963), .S0(d7_71__N_1531_adj_5700[38]), .S1(d7_71__N_1531_adj_5700[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1478_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1478_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1478_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_36 (.A0(d_d7_adj_5675[69]), .B0(d7_adj_5674[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[70]), .B1(d7_adj_5674[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16151), .COUT(n16152), .S0(n84_adj_5307), 
          .S1(n81_adj_5306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_32 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15750), .COUT(n15751), .S0(n96_adj_5043), .S1(n93_adj_5042));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_34 (.A0(d_d7_adj_5675[67]), .B0(d7_adj_5674[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[68]), .B1(d7_adj_5674[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16150), .COUT(n16151), .S0(n90_adj_5309), 
          .S1(n87_adj_5308));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_32 (.A0(d_d7_adj_5675[65]), .B0(d7_adj_5674[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[66]), .B1(d7_adj_5674[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16149), .COUT(n16150), .S0(n96_adj_5311), 
          .S1(n93_adj_5310));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_32.INJECT1_1 = "NO";
    CCU2C add_3644_15 (.A0(d_out_d_11__N_1875), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1875), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16399), .S0(n52), .S1(d_out_d_11__N_1878[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_15.INIT0 = 16'h666a;
    defparam add_3644_15.INIT1 = 16'h666a;
    defparam add_3644_15.INJECT1_0 = "NO";
    defparam add_3644_15.INJECT1_1 = "NO";
    CCU2C add_3644_13 (.A0(d_out_d_11__N_1876[17]), .B0(n51_adj_5553), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n48_adj_5552), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16398), .COUT(n16399), .S0(n58), 
          .S1(n55));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_13.INIT0 = 16'h9995;
    defparam add_3644_13.INIT1 = 16'h9995;
    defparam add_3644_13.INJECT1_0 = "NO";
    defparam add_3644_13.INJECT1_1 = "NO";
    CCU2C add_3644_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n57_adj_5555), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n54_adj_5554), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16397), .COUT(n16398), .S0(n64_adj_5378), 
          .S1(n61));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_11.INIT0 = 16'h6969;
    defparam add_3644_11.INIT1 = 16'h9995;
    defparam add_3644_11.INJECT1_0 = "NO";
    defparam add_3644_11.INJECT1_1 = "NO";
    CCU2C add_3644_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n63_adj_5557), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1876[17]), 
          .C1(n60_adj_5556), .D1(VCC_net), .CIN(n16396), .COUT(n16397), 
          .S0(n70), .S1(n67_adj_5379));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_9.INIT0 = 16'h6969;
    defparam add_3644_9.INIT1 = 16'h6969;
    defparam add_3644_9.INJECT1_0 = "NO";
    defparam add_3644_9.INJECT1_1 = "NO";
    CCU2C add_3644_7 (.A0(d_out_d_11__N_1876[17]), .B0(n17635), .C0(n69_adj_5559), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n66_adj_5558), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16395), .COUT(n16396), .S0(n76_adj_5380), 
          .S1(n73));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_7.INIT0 = 16'h6969;
    defparam add_3644_7.INIT1 = 16'h9995;
    defparam add_3644_7.INJECT1_0 = "NO";
    defparam add_3644_7.INJECT1_1 = "NO";
    CCU2C add_3644_5 (.A0(n75_adj_5561), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1876[17]), .C1(n72_adj_5560), 
          .D1(VCC_net), .CIN(n16394), .COUT(n16395), .S0(n82_adj_5382), 
          .S1(n79_adj_5381));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_5.INIT0 = 16'haaa0;
    defparam add_3644_5.INIT1 = 16'h9696;
    defparam add_3644_5.INJECT1_0 = "NO";
    defparam add_3644_5.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_30 (.A0(d_d7_adj_5675[63]), .B0(d7_adj_5674[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[64]), .B1(d7_adj_5674[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16148), .COUT(n16149), .S0(n102_adj_5313), 
          .S1(n99_adj_5312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_30.INJECT1_1 = "NO";
    LUT4 o_Rx_Byte_0__bdd_4_lut_3_lut (.A(o_Rx_Byte[3]), .B(o_Rx_Byte[2]), 
         .C(MYLED_0_6), .Z(n17522)) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_0__bdd_4_lut_3_lut.init = 16'h6f6f;
    CCU2C add_3644_3 (.A0(d_out_d_11__N_1876[17]), .B0(ISquare[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16393), .COUT(n16394), .S1(n85_adj_5383));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_3.INIT0 = 16'h666a;
    defparam add_3644_3.INIT1 = 16'h555f;
    defparam add_3644_3.INJECT1_0 = "NO";
    defparam add_3644_3.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_35 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15845), .COUT(n15846), .S0(n82), .S1(n79));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_35.INJECT1_1 = "NO";
    CCU2C add_3644_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16393));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3644_1.INIT0 = 16'h0000;
    defparam add_3644_1.INIT1 = 16'haaaf;
    defparam add_3644_1.INJECT1_0 = "NO";
    defparam add_3644_1.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_30 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15749), .COUT(n15750), .S0(n102_adj_5045), .S1(n99_adj_5044));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_14 (.A0(d_d9_adj_5679[11]), .B0(d9_adj_5678[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[12]), .B1(d9_adj_5678[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15558), .COUT(n15559));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_12 (.A0(d_d9_adj_5679[9]), .B0(d9_adj_5678[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[10]), .B1(d9_adj_5678[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15557), .COUT(n15558));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_10 (.A0(d_d9_adj_5679[7]), .B0(d9_adj_5678[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[8]), .B1(d9_adj_5678[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15556), .COUT(n15557));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_8 (.A0(d_d9_adj_5679[5]), .B0(d9_adj_5678[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[6]), .B1(d9_adj_5678[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15555), .COUT(n15556));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_6 (.A0(d_d9_adj_5679[3]), .B0(d9_adj_5678[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[4]), .B1(d9_adj_5678[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15554), .COUT(n15555));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_4 (.A0(d_d9_adj_5679[1]), .B0(d9_adj_5678[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[2]), .B1(d9_adj_5678[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15553), .COUT(n15554));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5679[0]), .B1(d9_adj_5678[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15553));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1595_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1595_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_37 (.A0(d3_adj_5669[70]), .B0(cout_adj_5136), 
          .C0(n81_adj_4564), .D0(d4_adj_5670[70]), .A1(d3_adj_5669[71]), 
          .B1(cout_adj_5136), .C1(n78_adj_4565), .D1(d4_adj_5670[71]), 
          .CIN(n15551), .S0(d4_71__N_634_adj_5686[70]), .S1(d4_71__N_634_adj_5686[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_35 (.A0(d3_adj_5669[68]), .B0(cout_adj_5136), 
          .C0(n87_adj_4562), .D0(d4_adj_5670[68]), .A1(d3_adj_5669[69]), 
          .B1(cout_adj_5136), .C1(n84_adj_4563), .D1(d4_adj_5670[69]), 
          .CIN(n15550), .COUT(n15551), .S0(d4_71__N_634_adj_5686[68]), 
          .S1(d4_71__N_634_adj_5686[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_33 (.A0(d3_adj_5669[66]), .B0(cout_adj_5136), 
          .C0(n93_adj_4560), .D0(d4_adj_5670[66]), .A1(d3_adj_5669[67]), 
          .B1(cout_adj_5136), .C1(n90_adj_4561), .D1(d4_adj_5670[67]), 
          .CIN(n15549), .COUT(n15550), .S0(d4_71__N_634_adj_5686[66]), 
          .S1(d4_71__N_634_adj_5686[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_31 (.A0(d3_adj_5669[64]), .B0(cout_adj_5136), 
          .C0(n99_adj_4558), .D0(d4_adj_5670[64]), .A1(d3_adj_5669[65]), 
          .B1(cout_adj_5136), .C1(n96_adj_4559), .D1(d4_adj_5670[65]), 
          .CIN(n15548), .COUT(n15549), .S0(d4_71__N_634_adj_5686[64]), 
          .S1(d4_71__N_634_adj_5686[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_29 (.A0(d3_adj_5669[62]), .B0(cout_adj_5136), 
          .C0(n105_adj_4556), .D0(d4_adj_5670[62]), .A1(d3_adj_5669[63]), 
          .B1(cout_adj_5136), .C1(n102_adj_4557), .D1(d4_adj_5670[63]), 
          .CIN(n15547), .COUT(n15548), .S0(d4_71__N_634_adj_5686[62]), 
          .S1(d4_71__N_634_adj_5686[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_27 (.A0(d3_adj_5669[60]), .B0(cout_adj_5136), 
          .C0(n111_adj_4554), .D0(d4_adj_5670[60]), .A1(d3_adj_5669[61]), 
          .B1(cout_adj_5136), .C1(n108_adj_4555), .D1(d4_adj_5670[61]), 
          .CIN(n15546), .COUT(n15547), .S0(d4_71__N_634_adj_5686[60]), 
          .S1(d4_71__N_634_adj_5686[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_25 (.A0(d3_adj_5669[58]), .B0(cout_adj_5136), 
          .C0(n117_adj_4552), .D0(d4_adj_5670[58]), .A1(d3_adj_5669[59]), 
          .B1(cout_adj_5136), .C1(n114_adj_4553), .D1(d4_adj_5670[59]), 
          .CIN(n15545), .COUT(n15546), .S0(d4_71__N_634_adj_5686[58]), 
          .S1(d4_71__N_634_adj_5686[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_23 (.A0(d3_adj_5669[56]), .B0(cout_adj_5136), 
          .C0(n123_adj_4550), .D0(d4_adj_5670[56]), .A1(d3_adj_5669[57]), 
          .B1(cout_adj_5136), .C1(n120_adj_4551), .D1(d4_adj_5670[57]), 
          .CIN(n15544), .COUT(n15545), .S0(d4_71__N_634_adj_5686[56]), 
          .S1(d4_71__N_634_adj_5686[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_21 (.A0(d3_adj_5669[54]), .B0(cout_adj_5136), 
          .C0(n129_adj_4548), .D0(d4_adj_5670[54]), .A1(d3_adj_5669[55]), 
          .B1(cout_adj_5136), .C1(n126_adj_4549), .D1(d4_adj_5670[55]), 
          .CIN(n15543), .COUT(n15544), .S0(d4_71__N_634_adj_5686[54]), 
          .S1(d4_71__N_634_adj_5686[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_19 (.A0(d3_adj_5669[52]), .B0(cout_adj_5136), 
          .C0(n135_adj_4546), .D0(d4_adj_5670[52]), .A1(d3_adj_5669[53]), 
          .B1(cout_adj_5136), .C1(n132_adj_4547), .D1(d4_adj_5670[53]), 
          .CIN(n15542), .COUT(n15543), .S0(d4_71__N_634_adj_5686[52]), 
          .S1(d4_71__N_634_adj_5686[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_17 (.A0(d3_adj_5669[50]), .B0(cout_adj_5136), 
          .C0(n141_adj_4544), .D0(d4_adj_5670[50]), .A1(d3_adj_5669[51]), 
          .B1(cout_adj_5136), .C1(n138_adj_4545), .D1(d4_adj_5670[51]), 
          .CIN(n15541), .COUT(n15542), .S0(d4_71__N_634_adj_5686[50]), 
          .S1(d4_71__N_634_adj_5686[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_15 (.A0(d3_adj_5669[48]), .B0(cout_adj_5136), 
          .C0(n147_adj_4542), .D0(d4_adj_5670[48]), .A1(d3_adj_5669[49]), 
          .B1(cout_adj_5136), .C1(n144_adj_4543), .D1(d4_adj_5670[49]), 
          .CIN(n15540), .COUT(n15541), .S0(d4_71__N_634_adj_5686[48]), 
          .S1(d4_71__N_634_adj_5686[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_13 (.A0(d3_adj_5669[46]), .B0(cout_adj_5136), 
          .C0(n153_adj_4540), .D0(d4_adj_5670[46]), .A1(d3_adj_5669[47]), 
          .B1(cout_adj_5136), .C1(n150_adj_4541), .D1(d4_adj_5670[47]), 
          .CIN(n15539), .COUT(n15540), .S0(d4_71__N_634_adj_5686[46]), 
          .S1(d4_71__N_634_adj_5686[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_11 (.A0(d3_adj_5669[44]), .B0(cout_adj_5136), 
          .C0(n159_adj_3855), .D0(d4_adj_5670[44]), .A1(d3_adj_5669[45]), 
          .B1(cout_adj_5136), .C1(n156_adj_4520), .D1(d4_adj_5670[45]), 
          .CIN(n15538), .COUT(n15539), .S0(d4_71__N_634_adj_5686[44]), 
          .S1(d4_71__N_634_adj_5686[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_9 (.A0(d3_adj_5669[42]), .B0(cout_adj_5136), 
          .C0(n165), .D0(d4_adj_5670[42]), .A1(d3_adj_5669[43]), .B1(cout_adj_5136), 
          .C1(n162_adj_3854), .D1(d4_adj_5670[43]), .CIN(n15537), .COUT(n15538), 
          .S0(d4_71__N_634_adj_5686[42]), .S1(d4_71__N_634_adj_5686[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_7 (.A0(d3_adj_5669[40]), .B0(cout_adj_5136), 
          .C0(n171), .D0(d4_adj_5670[40]), .A1(d3_adj_5669[41]), .B1(cout_adj_5136), 
          .C1(n168), .D1(d4_adj_5670[41]), .CIN(n15536), .COUT(n15537), 
          .S0(d4_71__N_634_adj_5686[40]), .S1(d4_71__N_634_adj_5686[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_5 (.A0(d3_adj_5669[38]), .B0(cout_adj_5136), 
          .C0(n177), .D0(d4_adj_5670[38]), .A1(d3_adj_5669[39]), .B1(cout_adj_5136), 
          .C1(n174), .D1(d4_adj_5670[39]), .CIN(n15535), .COUT(n15536), 
          .S0(d4_71__N_634_adj_5686[38]), .S1(d4_71__N_634_adj_5686[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_3 (.A0(d3_adj_5669[36]), .B0(cout_adj_5136), 
          .C0(n183_adj_4539), .D0(d4_adj_5670[36]), .A1(d3_adj_5669[37]), 
          .B1(cout_adj_5136), .C1(n180), .D1(d4_adj_5670[37]), .CIN(n15534), 
          .COUT(n15535), .S0(d4_71__N_634_adj_5686[36]), .S1(d4_71__N_634_adj_5686[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1493_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1493_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5136), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15534));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1493_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1493_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1493_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_13 (.A0(LOCosine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15530), .S0(MixerOutCos_11__N_250[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1457_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1457_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_11 (.A0(LOCosine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15529), .COUT(n15530), .S0(MixerOutCos_11__N_250[9]), 
          .S1(MixerOutCos_11__N_250[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1457_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1457_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_9 (.A0(LOCosine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15528), .COUT(n15529), .S0(MixerOutCos_11__N_250[7]), 
          .S1(MixerOutCos_11__N_250[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1457_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1457_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_7 (.A0(LOCosine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15527), .COUT(n15528), .S0(MixerOutCos_11__N_250[5]), 
          .S1(MixerOutCos_11__N_250[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1457_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1457_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_5 (.A0(LOCosine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15526), .COUT(n15527), .S0(MixerOutCos_11__N_250[3]), 
          .S1(MixerOutCos_11__N_250[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1457_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1457_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_3 (.A0(LOCosine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15525), .COUT(n15526), .S0(MixerOutCos_11__N_250[1]), 
          .S1(MixerOutCos_11__N_250[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1457_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1457_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15525), .S1(MixerOutCos_11__N_250[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(42[26:33])
    defparam _add_1_1457_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1457_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1457_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_63 (.A0(phase_inc_carrGen[62]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15523), .S0(n133), .S1(n130));
    defparam _add_1_1412_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_61 (.A0(phase_inc_carrGen[60]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15522), .COUT(n15523), .S0(n139), 
          .S1(n136));
    defparam _add_1_1412_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_59 (.A0(phase_inc_carrGen[58]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15521), .COUT(n15522), .S0(n145), 
          .S1(n142));
    defparam _add_1_1412_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_57 (.A0(phase_inc_carrGen[56]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15520), .COUT(n15521), .S0(n151), 
          .S1(n148));
    defparam _add_1_1412_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_55 (.A0(phase_inc_carrGen[54]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15519), .COUT(n15520), .S0(n157), 
          .S1(n154));
    defparam _add_1_1412_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_53 (.A0(phase_inc_carrGen[52]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15518), .COUT(n15519), .S0(n163), 
          .S1(n160));
    defparam _add_1_1412_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_51 (.A0(phase_inc_carrGen[50]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15517), .COUT(n15518), .S0(n169), 
          .S1(n166));
    defparam _add_1_1412_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_49 (.A0(phase_inc_carrGen[48]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15516), .COUT(n15517), .S0(n175), 
          .S1(n172));
    defparam _add_1_1412_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_47 (.A0(phase_inc_carrGen[46]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15515), .COUT(n15516), .S0(n181), 
          .S1(n178));
    defparam _add_1_1412_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_45 (.A0(phase_inc_carrGen[44]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15514), .COUT(n15515), .S0(n187), 
          .S1(n184));
    defparam _add_1_1412_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_43 (.A0(phase_inc_carrGen[42]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15513), .COUT(n15514), .S0(n193), 
          .S1(n190));
    defparam _add_1_1412_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_41 (.A0(phase_inc_carrGen[40]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15512), .COUT(n15513), .S0(n199), 
          .S1(n196));
    defparam _add_1_1412_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_39 (.A0(phase_inc_carrGen[38]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15511), .COUT(n15512), .S0(n205), 
          .S1(n202));
    defparam _add_1_1412_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_37 (.A0(phase_inc_carrGen[36]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15510), .COUT(n15511), .S0(n211), 
          .S1(n208));
    defparam _add_1_1412_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_35 (.A0(phase_inc_carrGen[34]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15509), .COUT(n15510), .S0(n217), 
          .S1(n214));
    defparam _add_1_1412_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_33 (.A0(phase_inc_carrGen[32]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15508), .COUT(n15509), .S0(n223), 
          .S1(n220));
    defparam _add_1_1412_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_31 (.A0(phase_inc_carrGen[30]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15507), .COUT(n15508), .S0(n229), 
          .S1(n226));
    defparam _add_1_1412_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_29 (.A0(phase_inc_carrGen[28]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15506), .COUT(n15507), .S0(n235), 
          .S1(n232));
    defparam _add_1_1412_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_27 (.A0(phase_inc_carrGen[26]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15505), .COUT(n15506), .S0(n241), 
          .S1(n238));
    defparam _add_1_1412_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_25 (.A0(phase_inc_carrGen[24]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15504), .COUT(n15505), .S0(n247), 
          .S1(n244));
    defparam _add_1_1412_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_23 (.A0(phase_inc_carrGen[22]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15503), .COUT(n15504), .S0(n253), 
          .S1(n250));
    defparam _add_1_1412_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_21 (.A0(phase_inc_carrGen[20]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15502), .COUT(n15503), .S0(n259), 
          .S1(n256));
    defparam _add_1_1412_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_19 (.A0(phase_inc_carrGen[18]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15501), .COUT(n15502), .S0(n265), 
          .S1(n262));
    defparam _add_1_1412_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_17 (.A0(phase_inc_carrGen[16]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15500), .COUT(n15501), .S0(n271), 
          .S1(n268));
    defparam _add_1_1412_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_15 (.A0(phase_inc_carrGen[14]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15499), .COUT(n15500), .S0(n277), 
          .S1(n274));
    defparam _add_1_1412_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_13 (.A0(phase_inc_carrGen[12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15498), .COUT(n15499), .S0(n283), 
          .S1(n280));
    defparam _add_1_1412_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_1412_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_11 (.A0(phase_inc_carrGen[10]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15497), .COUT(n15498), .S0(n289), 
          .S1(n286));
    defparam _add_1_1412_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_9 (.A0(phase_inc_carrGen[8]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15496), .COUT(n15497), .S0(n295), 
          .S1(n292));
    defparam _add_1_1412_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_9.INJECT1_1 = "NO";
    CCU2C add_3637_19 (.A0(d_out_d_11__N_1882[17]), .B0(n48_adj_5490), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n45_adj_5489), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16387), .S0(n45_adj_5473), 
          .S1(d_out_d_11__N_1884[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_19.INIT0 = 16'h9995;
    defparam add_3637_19.INIT1 = 16'h9995;
    defparam add_3637_19.INJECT1_0 = "NO";
    defparam add_3637_19.INJECT1_1 = "NO";
    CCU2C add_3637_17 (.A0(d_out_d_11__N_1882[17]), .B0(n54_adj_5492), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n51_adj_5491), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16386), .COUT(n16387), .S0(n51_adj_5475), 
          .S1(n48_adj_5474));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_17.INIT0 = 16'h9995;
    defparam add_3637_17.INIT1 = 16'h9995;
    defparam add_3637_17.INJECT1_0 = "NO";
    defparam add_3637_17.INJECT1_1 = "NO";
    CCU2C add_3637_15 (.A0(d_out_d_11__N_1882[17]), .B0(n60_adj_5494), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n57_adj_5493), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16385), .COUT(n16386), .S0(n57_adj_5477), 
          .S1(n54_adj_5476));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_15.INIT0 = 16'h9995;
    defparam add_3637_15.INIT1 = 16'h9995;
    defparam add_3637_15.INJECT1_0 = "NO";
    defparam add_3637_15.INJECT1_1 = "NO";
    CCU2C add_3637_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1882[17]), .C0(n66_adj_5496), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n63_adj_5495), .D1(VCC_net), .CIN(n16384), .COUT(n16385), 
          .S0(n63_adj_5479), .S1(n60_adj_5478));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_13.INIT0 = 16'h6969;
    defparam add_3637_13.INIT1 = 16'h6969;
    defparam add_3637_13.INJECT1_0 = "NO";
    defparam add_3637_13.INJECT1_1 = "NO";
    CCU2C add_3637_11 (.A0(d_out_d_11__N_1882[17]), .B0(n72_adj_5498), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n69_adj_5497), .D1(VCC_net), .CIN(n16383), .COUT(n16384), 
          .S0(n69_adj_5481), .S1(n66_adj_5480));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_11.INIT0 = 16'h9995;
    defparam add_3637_11.INIT1 = 16'h6969;
    defparam add_3637_11.INJECT1_0 = "NO";
    defparam add_3637_11.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_28 (.A0(d_d7_adj_5675[61]), .B0(d7_adj_5674[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[62]), .B1(d7_adj_5674[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16147), .COUT(n16148), .S0(n108_adj_5315), 
          .S1(n105_adj_5314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_26 (.A0(d_d7_adj_5675[59]), .B0(d7_adj_5674[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[60]), .B1(d7_adj_5674[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16146), .COUT(n16147), .S0(n114_adj_5317), 
          .S1(n111_adj_5316));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_24 (.A0(d_d7_adj_5675[57]), .B0(d7_adj_5674[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[58]), .B1(d7_adj_5674[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16145), .COUT(n16146), .S0(n120_adj_5319), 
          .S1(n117_adj_5318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_22 (.A0(d_d7_adj_5675[55]), .B0(d7_adj_5674[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[56]), .B1(d7_adj_5674[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16144), .COUT(n16145), .S0(n126_adj_5321), 
          .S1(n123_adj_5320));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_20 (.A0(d_d7_adj_5675[53]), .B0(d7_adj_5674[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[54]), .B1(d7_adj_5674[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16143), .COUT(n16144), .S0(n132_adj_5323), 
          .S1(n129_adj_5322));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_18 (.A0(d_d7_adj_5675[51]), .B0(d7_adj_5674[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[52]), .B1(d7_adj_5674[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16142), .COUT(n16143), .S0(n138_adj_5325), 
          .S1(n135_adj_5324));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_16 (.A0(d_d7_adj_5675[49]), .B0(d7_adj_5674[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[50]), .B1(d7_adj_5674[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16141), .COUT(n16142), .S0(n144_adj_5327), 
          .S1(n141_adj_5326));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_14 (.A0(d_d7_adj_5675[47]), .B0(d7_adj_5674[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[48]), .B1(d7_adj_5674[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16140), .COUT(n16141), .S0(n150_adj_5329), 
          .S1(n147_adj_5328));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_12 (.A0(d_d7_adj_5675[45]), .B0(d7_adj_5674[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[46]), .B1(d7_adj_5674[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16139), .COUT(n16140), .S0(n156_adj_5331), 
          .S1(n153_adj_5330));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_12.INJECT1_1 = "NO";
    CCU2C add_3637_9 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n78_adj_5500), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(n17635), .C1(n75_adj_5499), .D1(VCC_net), .CIN(n16382), 
          .COUT(n16383), .S0(n75_adj_5483), .S1(n72_adj_5482));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_9.INIT0 = 16'h9696;
    defparam add_3637_9.INIT1 = 16'h6969;
    defparam add_3637_9.INJECT1_0 = "NO";
    defparam add_3637_9.INJECT1_1 = "NO";
    CCU2C add_3637_7 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n84_adj_5502), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(n81_adj_5501), .D1(VCC_net), 
          .CIN(n16381), .COUT(n16382), .S0(n81_adj_5485), .S1(n78_adj_5484));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_7.INIT0 = 16'h9696;
    defparam add_3637_7.INIT1 = 16'h9696;
    defparam add_3637_7.INJECT1_0 = "NO";
    defparam add_3637_7.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_25 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n117_adj_5103), .D0(d1[58]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n114_adj_5102), .D1(d1[59]), .CIN(n15861), .COUT(n15862), 
          .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_25.INJECT1_1 = "NO";
    CCU2C add_3637_5 (.A0(n90_adj_5504), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1882[17]), .C1(n87_adj_5503), 
          .D1(VCC_net), .CIN(n16380), .COUT(n16381), .S0(n87_adj_5487), 
          .S1(n84_adj_5486));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_5.INIT0 = 16'haaa0;
    defparam add_3637_5.INIT1 = 16'h9696;
    defparam add_3637_5.INJECT1_0 = "NO";
    defparam add_3637_5.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_13 (.A0(d6[46]), .B0(cout_adj_5341), .C0(n153_adj_4950), 
          .D0(n27_adj_4708), .A1(d6[47]), .B1(cout_adj_5341), .C1(n150_adj_4949), 
          .D1(n26_adj_4709), .CIN(n16007), .COUT(n16008), .S0(d7_71__N_1531[46]), 
          .S1(d7_71__N_1531[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_13.INJECT1_1 = "NO";
    CCU2C add_3637_3 (.A0(d_out_d_11__N_1882[17]), .B0(ISquare[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16379), .COUT(n16380), .S1(n90_adj_5488));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_3.INIT0 = 16'h666a;
    defparam add_3637_3.INIT1 = 16'h555f;
    defparam add_3637_3.INJECT1_0 = "NO";
    defparam add_3637_3.INJECT1_1 = "NO";
    CCU2C add_3637_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16379));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3637_1.INIT0 = 16'h0000;
    defparam add_3637_1.INIT1 = 16'haaaf;
    defparam add_3637_1.INJECT1_0 = "NO";
    defparam add_3637_1.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_6 (.A0(MultResult2[4]), .B0(MultResult1[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[5]), .B1(MultResult1[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15796), .COUT(n15797), .S0(n114_adj_5174), 
          .S1(n111_adj_5173));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_6.INIT0 = 16'h666a;
    defparam ISquare_add_4_6.INIT1 = 16'h666a;
    defparam ISquare_add_4_6.INJECT1_0 = "NO";
    defparam ISquare_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_10 (.A0(d_d7_adj_5675[43]), .B0(d7_adj_5674[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[44]), .B1(d7_adj_5674[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16138), .COUT(n16139), .S0(n162_adj_5333), 
          .S1(n159_adj_5332));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_10.INJECT1_1 = "NO";
    CCU2C add_3639_17 (.A0(ISquare[31]), .B0(n913), .C0(GND_net), .D0(VCC_net), 
          .A1(n912), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16373), 
          .S1(d_out_d_11__N_2353[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_17.INIT0 = 16'h666a;
    defparam add_3639_17.INIT1 = 16'haaa0;
    defparam add_3639_17.INJECT1_0 = "NO";
    defparam add_3639_17.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_4 (.A0(MultResult2[2]), .B0(MultResult1[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[3]), .B1(MultResult1[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15795), .COUT(n15796), .S0(n120_adj_5176), 
          .S1(n117_adj_5175));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_4.INIT0 = 16'h666a;
    defparam ISquare_add_4_4.INIT1 = 16'h666a;
    defparam ISquare_add_4_4.INJECT1_0 = "NO";
    defparam ISquare_add_4_4.INJECT1_1 = "NO";
    CCU2C add_3639_15 (.A0(ISquare[31]), .B0(n915), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n914), .C1(GND_net), .D1(VCC_net), .CIN(n16372), 
          .COUT(n16373));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_15.INIT0 = 16'h666a;
    defparam add_3639_15.INIT1 = 16'h666a;
    defparam add_3639_15.INJECT1_0 = "NO";
    defparam add_3639_15.INJECT1_1 = "NO";
    CCU2C add_3639_13 (.A0(n917), .B0(n14874), .C0(n209), .D0(ISquare[31]), 
          .A1(n916), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16371), 
          .COUT(n16372));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_13.INIT0 = 16'h556a;
    defparam add_3639_13.INIT1 = 16'haaa0;
    defparam add_3639_13.INJECT1_0 = "NO";
    defparam add_3639_13.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_33 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15844), .COUT(n15845), .S0(n88), .S1(n85));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_33.INJECT1_1 = "NO";
    CCU2C add_3639_11 (.A0(d_out_d_11__N_1876[17]), .B0(n919), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n918), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16370), .COUT(n16371));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_11.INIT0 = 16'h9995;
    defparam add_3639_11.INIT1 = 16'h9995;
    defparam add_3639_11.INJECT1_0 = "NO";
    defparam add_3639_11.INJECT1_1 = "NO";
    CCU2C add_3639_9 (.A0(d_out_d_11__N_1880[17]), .B0(n921), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n920), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16369), .COUT(n16370));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_9.INIT0 = 16'h9995;
    defparam add_3639_9.INIT1 = 16'h9995;
    defparam add_3639_9.INJECT1_0 = "NO";
    defparam add_3639_9.INJECT1_1 = "NO";
    CCU2C add_3639_7 (.A0(d_out_d_11__N_1884[17]), .B0(n923), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n922), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16368), .COUT(n16369));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_7.INIT0 = 16'h9995;
    defparam add_3639_7.INIT1 = 16'h9995;
    defparam add_3639_7.INJECT1_0 = "NO";
    defparam add_3639_7.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_2 (.A0(MultResult2[0]), .B0(MultResult1[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[1]), .B1(MultResult1[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15795), .S1(n123_adj_5177));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_2.INIT0 = 16'h0008;
    defparam ISquare_add_4_2.INIT1 = 16'h666a;
    defparam ISquare_add_4_2.INJECT1_0 = "NO";
    defparam ISquare_add_4_2.INJECT1_1 = "NO";
    CCU2C add_3639_5 (.A0(d_out_d_11__N_1888[17]), .B0(n925), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n924), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16367), .COUT(n16368));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_5.INIT0 = 16'h9995;
    defparam add_3639_5.INIT1 = 16'h9995;
    defparam add_3639_5.INJECT1_0 = "NO";
    defparam add_3639_5.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_31 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15843), .COUT(n15844), .S0(n94), .S1(n91));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1484_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_31.INJECT1_1 = "NO";
    CCU2C add_3639_3 (.A0(d_out_d_11__N_1892[17]), .B0(n927), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n926), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16366), .COUT(n16367));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_3.INIT0 = 16'h9995;
    defparam add_3639_3.INIT1 = 16'h9995;
    defparam add_3639_3.INJECT1_0 = "NO";
    defparam add_3639_3.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_28 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15748), .COUT(n15749), .S0(n108_adj_5047), .S1(n105_adj_5046));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_28.INJECT1_1 = "NO";
    LUT4 mux_325_i4_3_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(n2636), .C(n310), 
         .D(n17629), .Z(n2367)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam mux_325_i4_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2C _add_1_1583_add_4_26 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15747), .COUT(n15748), .S0(n114_adj_5049), .S1(n111_adj_5048));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_24 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15746), .COUT(n15747), .S0(n120_adj_5051), .S1(n117_adj_5050));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_7 (.A0(phase_inc_carrGen[6]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15495), .COUT(n15496), .S0(n301), 
          .S1(n298));
    defparam _add_1_1412_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_5 (.A0(phase_inc_carrGen[4]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15494), .COUT(n15495), .S0(n307), 
          .S1(n304));
    defparam _add_1_1412_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_3 (.A0(phase_inc_carrGen[2]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[3]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15493), .COUT(n15494), .S0(n313), 
          .S1(n310));
    defparam _add_1_1412_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1412_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1412_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15493), .S1(n316));
    defparam _add_1_1412_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1412_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1412_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_38 (.A0(d_d_tmp_adj_5666[35]), .B0(d_tmp_adj_5665[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15492), .S0(d6_71__N_1459_adj_5699[35]), 
          .S1(cout_adj_5420));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1613_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_36 (.A0(d_d_tmp_adj_5666[33]), .B0(d_tmp_adj_5665[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[34]), .B1(d_tmp_adj_5665[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15491), .COUT(n15492), .S0(d6_71__N_1459_adj_5699[33]), 
          .S1(d6_71__N_1459_adj_5699[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_34 (.A0(d_d_tmp_adj_5666[31]), .B0(d_tmp_adj_5665[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[32]), .B1(d_tmp_adj_5665[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15490), .COUT(n15491), .S0(d6_71__N_1459_adj_5699[31]), 
          .S1(d6_71__N_1459_adj_5699[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_32 (.A0(d_d_tmp_adj_5666[29]), .B0(d_tmp_adj_5665[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[30]), .B1(d_tmp_adj_5665[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15489), .COUT(n15490), .S0(d6_71__N_1459_adj_5699[29]), 
          .S1(d6_71__N_1459_adj_5699[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_30 (.A0(d_d_tmp_adj_5666[27]), .B0(d_tmp_adj_5665[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[28]), .B1(d_tmp_adj_5665[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15488), .COUT(n15489), .S0(d6_71__N_1459_adj_5699[27]), 
          .S1(d6_71__N_1459_adj_5699[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_28 (.A0(d_d_tmp_adj_5666[25]), .B0(d_tmp_adj_5665[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[26]), .B1(d_tmp_adj_5665[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15487), .COUT(n15488), .S0(d6_71__N_1459_adj_5699[25]), 
          .S1(d6_71__N_1459_adj_5699[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_26 (.A0(d_d_tmp_adj_5666[23]), .B0(d_tmp_adj_5665[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[24]), .B1(d_tmp_adj_5665[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15486), .COUT(n15487), .S0(d6_71__N_1459_adj_5699[23]), 
          .S1(d6_71__N_1459_adj_5699[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_24 (.A0(d_d_tmp_adj_5666[21]), .B0(d_tmp_adj_5665[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[22]), .B1(d_tmp_adj_5665[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15485), .COUT(n15486), .S0(d6_71__N_1459_adj_5699[21]), 
          .S1(d6_71__N_1459_adj_5699[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_22 (.A0(d_d_tmp_adj_5666[19]), .B0(d_tmp_adj_5665[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[20]), .B1(d_tmp_adj_5665[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15484), .COUT(n15485), .S0(d6_71__N_1459_adj_5699[19]), 
          .S1(d6_71__N_1459_adj_5699[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_20 (.A0(d_d_tmp_adj_5666[17]), .B0(d_tmp_adj_5665[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[18]), .B1(d_tmp_adj_5665[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15483), .COUT(n15484), .S0(d6_71__N_1459_adj_5699[17]), 
          .S1(d6_71__N_1459_adj_5699[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_18 (.A0(d_d_tmp_adj_5666[15]), .B0(d_tmp_adj_5665[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[16]), .B1(d_tmp_adj_5665[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15482), .COUT(n15483), .S0(d6_71__N_1459_adj_5699[15]), 
          .S1(d6_71__N_1459_adj_5699[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_16 (.A0(d_d_tmp_adj_5666[13]), .B0(d_tmp_adj_5665[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[14]), .B1(d_tmp_adj_5665[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15481), .COUT(n15482), .S0(d6_71__N_1459_adj_5699[13]), 
          .S1(d6_71__N_1459_adj_5699[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_14 (.A0(d_d_tmp_adj_5666[11]), .B0(d_tmp_adj_5665[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[12]), .B1(d_tmp_adj_5665[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15480), .COUT(n15481), .S0(d6_71__N_1459_adj_5699[11]), 
          .S1(d6_71__N_1459_adj_5699[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_12 (.A0(d_d_tmp_adj_5666[9]), .B0(d_tmp_adj_5665[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[10]), .B1(d_tmp_adj_5665[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15479), .COUT(n15480), .S0(d6_71__N_1459_adj_5699[9]), 
          .S1(d6_71__N_1459_adj_5699[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_10 (.A0(d_d_tmp_adj_5666[7]), .B0(d_tmp_adj_5665[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[8]), .B1(d_tmp_adj_5665[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15478), .COUT(n15479), .S0(d6_71__N_1459_adj_5699[7]), 
          .S1(d6_71__N_1459_adj_5699[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_8 (.A0(d_d_tmp_adj_5666[5]), .B0(d_tmp_adj_5665[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[6]), .B1(d_tmp_adj_5665[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15477), .COUT(n15478), .S0(d6_71__N_1459_adj_5699[5]), 
          .S1(d6_71__N_1459_adj_5699[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_6 (.A0(d_d_tmp_adj_5666[3]), .B0(d_tmp_adj_5665[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[4]), .B1(d_tmp_adj_5665[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15476), .COUT(n15477), .S0(d6_71__N_1459_adj_5699[3]), 
          .S1(d6_71__N_1459_adj_5699[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_4 (.A0(d_d_tmp_adj_5666[1]), .B0(d_tmp_adj_5665[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[2]), .B1(d_tmp_adj_5665[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15475), .COUT(n15476), .S0(d6_71__N_1459_adj_5699[1]), 
          .S1(d6_71__N_1459_adj_5699[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1613_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1613_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5666[0]), .B1(d_tmp_adj_5665[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15475), .S1(d6_71__N_1459_adj_5699[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1613_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1613_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1613_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1613_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_37 (.A0(d2_adj_5668[70]), .B0(cout_adj_5135), 
          .C0(n81_adj_4839), .D0(d3_adj_5669[70]), .A1(d2_adj_5668[71]), 
          .B1(cout_adj_5135), .C1(n78_adj_4838), .D1(d3_adj_5669[71]), 
          .CIN(n15473), .S0(d3_71__N_562_adj_5685[70]), .S1(d3_71__N_562_adj_5685[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_35 (.A0(d2_adj_5668[68]), .B0(cout_adj_5135), 
          .C0(n87_adj_4841), .D0(d3_adj_5669[68]), .A1(d2_adj_5668[69]), 
          .B1(cout_adj_5135), .C1(n84_adj_4840), .D1(d3_adj_5669[69]), 
          .CIN(n15472), .COUT(n15473), .S0(d3_71__N_562_adj_5685[68]), 
          .S1(d3_71__N_562_adj_5685[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_33 (.A0(d2_adj_5668[66]), .B0(cout_adj_5135), 
          .C0(n93_adj_4843), .D0(d3_adj_5669[66]), .A1(d2_adj_5668[67]), 
          .B1(cout_adj_5135), .C1(n90_adj_4842), .D1(d3_adj_5669[67]), 
          .CIN(n15471), .COUT(n15472), .S0(d3_71__N_562_adj_5685[66]), 
          .S1(d3_71__N_562_adj_5685[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_31 (.A0(d2_adj_5668[64]), .B0(cout_adj_5135), 
          .C0(n99_adj_4845), .D0(d3_adj_5669[64]), .A1(d2_adj_5668[65]), 
          .B1(cout_adj_5135), .C1(n96_adj_4844), .D1(d3_adj_5669[65]), 
          .CIN(n15470), .COUT(n15471), .S0(d3_71__N_562_adj_5685[64]), 
          .S1(d3_71__N_562_adj_5685[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_29 (.A0(d2_adj_5668[62]), .B0(cout_adj_5135), 
          .C0(n105_adj_4847), .D0(d3_adj_5669[62]), .A1(d2_adj_5668[63]), 
          .B1(cout_adj_5135), .C1(n102_adj_4846), .D1(d3_adj_5669[63]), 
          .CIN(n15469), .COUT(n15470), .S0(d3_71__N_562_adj_5685[62]), 
          .S1(d3_71__N_562_adj_5685[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_27 (.A0(d2_adj_5668[60]), .B0(cout_adj_5135), 
          .C0(n111_adj_4849), .D0(d3_adj_5669[60]), .A1(d2_adj_5668[61]), 
          .B1(cout_adj_5135), .C1(n108_adj_4848), .D1(d3_adj_5669[61]), 
          .CIN(n15468), .COUT(n15469), .S0(d3_71__N_562_adj_5685[60]), 
          .S1(d3_71__N_562_adj_5685[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_25 (.A0(d2_adj_5668[58]), .B0(cout_adj_5135), 
          .C0(n117_adj_4851), .D0(d3_adj_5669[58]), .A1(d2_adj_5668[59]), 
          .B1(cout_adj_5135), .C1(n114_adj_4850), .D1(d3_adj_5669[59]), 
          .CIN(n15467), .COUT(n15468), .S0(d3_71__N_562_adj_5685[58]), 
          .S1(d3_71__N_562_adj_5685[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_23 (.A0(d2_adj_5668[56]), .B0(cout_adj_5135), 
          .C0(n123_adj_4853), .D0(d3_adj_5669[56]), .A1(d2_adj_5668[57]), 
          .B1(cout_adj_5135), .C1(n120_adj_4852), .D1(d3_adj_5669[57]), 
          .CIN(n15466), .COUT(n15467), .S0(d3_71__N_562_adj_5685[56]), 
          .S1(d3_71__N_562_adj_5685[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_21 (.A0(d2_adj_5668[54]), .B0(cout_adj_5135), 
          .C0(n129_adj_4855), .D0(d3_adj_5669[54]), .A1(d2_adj_5668[55]), 
          .B1(cout_adj_5135), .C1(n126_adj_4854), .D1(d3_adj_5669[55]), 
          .CIN(n15465), .COUT(n15466), .S0(d3_71__N_562_adj_5685[54]), 
          .S1(d3_71__N_562_adj_5685[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_19 (.A0(d2_adj_5668[52]), .B0(cout_adj_5135), 
          .C0(n135_adj_4857), .D0(d3_adj_5669[52]), .A1(d2_adj_5668[53]), 
          .B1(cout_adj_5135), .C1(n132_adj_4856), .D1(d3_adj_5669[53]), 
          .CIN(n15464), .COUT(n15465), .S0(d3_71__N_562_adj_5685[52]), 
          .S1(d3_71__N_562_adj_5685[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_17 (.A0(d2_adj_5668[50]), .B0(cout_adj_5135), 
          .C0(n141_adj_4859), .D0(d3_adj_5669[50]), .A1(d2_adj_5668[51]), 
          .B1(cout_adj_5135), .C1(n138_adj_4858), .D1(d3_adj_5669[51]), 
          .CIN(n15463), .COUT(n15464), .S0(d3_71__N_562_adj_5685[50]), 
          .S1(d3_71__N_562_adj_5685[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_15 (.A0(d2_adj_5668[48]), .B0(cout_adj_5135), 
          .C0(n147_adj_4861), .D0(d3_adj_5669[48]), .A1(d2_adj_5668[49]), 
          .B1(cout_adj_5135), .C1(n144_adj_4860), .D1(d3_adj_5669[49]), 
          .CIN(n15462), .COUT(n15463), .S0(d3_71__N_562_adj_5685[48]), 
          .S1(d3_71__N_562_adj_5685[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_13 (.A0(d2_adj_5668[46]), .B0(cout_adj_5135), 
          .C0(n153_adj_4863), .D0(d3_adj_5669[46]), .A1(d2_adj_5668[47]), 
          .B1(cout_adj_5135), .C1(n150_adj_4862), .D1(d3_adj_5669[47]), 
          .CIN(n15461), .COUT(n15462), .S0(d3_71__N_562_adj_5685[46]), 
          .S1(d3_71__N_562_adj_5685[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_11 (.A0(d2_adj_5668[44]), .B0(cout_adj_5135), 
          .C0(n159_adj_4865), .D0(d3_adj_5669[44]), .A1(d2_adj_5668[45]), 
          .B1(cout_adj_5135), .C1(n156_adj_4864), .D1(d3_adj_5669[45]), 
          .CIN(n15460), .COUT(n15461), .S0(d3_71__N_562_adj_5685[44]), 
          .S1(d3_71__N_562_adj_5685[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_9 (.A0(d2_adj_5668[42]), .B0(cout_adj_5135), 
          .C0(n165_adj_4867), .D0(d3_adj_5669[42]), .A1(d2_adj_5668[43]), 
          .B1(cout_adj_5135), .C1(n162_adj_4866), .D1(d3_adj_5669[43]), 
          .CIN(n15459), .COUT(n15460), .S0(d3_71__N_562_adj_5685[42]), 
          .S1(d3_71__N_562_adj_5685[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_7 (.A0(d2_adj_5668[40]), .B0(cout_adj_5135), 
          .C0(n171_adj_4869), .D0(d3_adj_5669[40]), .A1(d2_adj_5668[41]), 
          .B1(cout_adj_5135), .C1(n168_adj_4868), .D1(d3_adj_5669[41]), 
          .CIN(n15458), .COUT(n15459), .S0(d3_71__N_562_adj_5685[40]), 
          .S1(d3_71__N_562_adj_5685[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_5 (.A0(d2_adj_5668[38]), .B0(cout_adj_5135), 
          .C0(n177_adj_4871), .D0(d3_adj_5669[38]), .A1(d2_adj_5668[39]), 
          .B1(cout_adj_5135), .C1(n174_adj_4870), .D1(d3_adj_5669[39]), 
          .CIN(n15457), .COUT(n15458), .S0(d3_71__N_562_adj_5685[38]), 
          .S1(d3_71__N_562_adj_5685[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_3 (.A0(d2_adj_5668[36]), .B0(cout_adj_5135), 
          .C0(n183_adj_4873), .D0(d3_adj_5669[36]), .A1(d2_adj_5668[37]), 
          .B1(cout_adj_5135), .C1(n180_adj_4872), .D1(d3_adj_5669[37]), 
          .CIN(n15456), .COUT(n15457), .S0(d3_71__N_562_adj_5685[36]), 
          .S1(d3_71__N_562_adj_5685[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1496_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1496_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1496_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5135), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15456));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1496_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1496_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1496_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1496_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_38 (.A0(d_d6_adj_5673[35]), .B0(d6_adj_5672[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15452), .S0(d7_71__N_1531_adj_5700[35]), 
          .S1(cout_adj_5179));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1610_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_36 (.A0(d_d6_adj_5673[33]), .B0(d6_adj_5672[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[34]), .B1(d6_adj_5672[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15451), .COUT(n15452), .S0(d7_71__N_1531_adj_5700[33]), 
          .S1(d7_71__N_1531_adj_5700[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_34 (.A0(d_d6_adj_5673[31]), .B0(d6_adj_5672[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[32]), .B1(d6_adj_5672[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15450), .COUT(n15451), .S0(d7_71__N_1531_adj_5700[31]), 
          .S1(d7_71__N_1531_adj_5700[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_32 (.A0(d_d6_adj_5673[29]), .B0(d6_adj_5672[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[30]), .B1(d6_adj_5672[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15449), .COUT(n15450), .S0(d7_71__N_1531_adj_5700[29]), 
          .S1(d7_71__N_1531_adj_5700[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_30 (.A0(d_d6_adj_5673[27]), .B0(d6_adj_5672[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[28]), .B1(d6_adj_5672[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15448), .COUT(n15449), .S0(d7_71__N_1531_adj_5700[27]), 
          .S1(d7_71__N_1531_adj_5700[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_28 (.A0(d_d6_adj_5673[25]), .B0(d6_adj_5672[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[26]), .B1(d6_adj_5672[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15447), .COUT(n15448), .S0(d7_71__N_1531_adj_5700[25]), 
          .S1(d7_71__N_1531_adj_5700[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_26 (.A0(d_d6_adj_5673[23]), .B0(d6_adj_5672[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[24]), .B1(d6_adj_5672[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15446), .COUT(n15447), .S0(d7_71__N_1531_adj_5700[23]), 
          .S1(d7_71__N_1531_adj_5700[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_24 (.A0(d_d6_adj_5673[21]), .B0(d6_adj_5672[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[22]), .B1(d6_adj_5672[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15445), .COUT(n15446), .S0(d7_71__N_1531_adj_5700[21]), 
          .S1(d7_71__N_1531_adj_5700[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_22 (.A0(d_d6_adj_5673[19]), .B0(d6_adj_5672[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[20]), .B1(d6_adj_5672[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15444), .COUT(n15445), .S0(d7_71__N_1531_adj_5700[19]), 
          .S1(d7_71__N_1531_adj_5700[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_20 (.A0(d_d6_adj_5673[17]), .B0(d6_adj_5672[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[18]), .B1(d6_adj_5672[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15443), .COUT(n15444), .S0(d7_71__N_1531_adj_5700[17]), 
          .S1(d7_71__N_1531_adj_5700[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_18 (.A0(d_d6_adj_5673[15]), .B0(d6_adj_5672[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[16]), .B1(d6_adj_5672[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15442), .COUT(n15443), .S0(d7_71__N_1531_adj_5700[15]), 
          .S1(d7_71__N_1531_adj_5700[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_16 (.A0(d_d6_adj_5673[13]), .B0(d6_adj_5672[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[14]), .B1(d6_adj_5672[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15441), .COUT(n15442), .S0(d7_71__N_1531_adj_5700[13]), 
          .S1(d7_71__N_1531_adj_5700[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_14 (.A0(d_d6_adj_5673[11]), .B0(d6_adj_5672[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[12]), .B1(d6_adj_5672[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15440), .COUT(n15441), .S0(d7_71__N_1531_adj_5700[11]), 
          .S1(d7_71__N_1531_adj_5700[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_12 (.A0(d_d6_adj_5673[9]), .B0(d6_adj_5672[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[10]), .B1(d6_adj_5672[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15439), .COUT(n15440), .S0(d7_71__N_1531_adj_5700[9]), 
          .S1(d7_71__N_1531_adj_5700[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_10 (.A0(d_d6_adj_5673[7]), .B0(d6_adj_5672[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[8]), .B1(d6_adj_5672[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15438), .COUT(n15439), .S0(d7_71__N_1531_adj_5700[7]), 
          .S1(d7_71__N_1531_adj_5700[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_8 (.A0(d_d6_adj_5673[5]), .B0(d6_adj_5672[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[6]), .B1(d6_adj_5672[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15437), .COUT(n15438), .S0(d7_71__N_1531_adj_5700[5]), 
          .S1(d7_71__N_1531_adj_5700[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_6 (.A0(d_d6_adj_5673[3]), .B0(d6_adj_5672[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[4]), .B1(d6_adj_5672[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15436), .COUT(n15437), .S0(d7_71__N_1531_adj_5700[3]), 
          .S1(d7_71__N_1531_adj_5700[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_4 (.A0(d_d6_adj_5673[1]), .B0(d6_adj_5672[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5673[2]), .B1(d6_adj_5672[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15435), .COUT(n15436), .S0(d7_71__N_1531_adj_5700[1]), 
          .S1(d7_71__N_1531_adj_5700[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1610_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1610_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5673[0]), .B1(d6_adj_5672[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15435), .S1(d7_71__N_1531_adj_5700[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1610_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1610_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1610_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1610_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_37 (.A0(d1_adj_5667[70]), .B0(cout_adj_5134), 
          .C0(n81_adj_5563), .D0(d2_adj_5668[70]), .A1(d1_adj_5667[71]), 
          .B1(cout_adj_5134), .C1(n78_adj_5562), .D1(d2_adj_5668[71]), 
          .CIN(n15433), .S0(d2_71__N_490_adj_5684[70]), .S1(d2_71__N_490_adj_5684[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_35 (.A0(d1_adj_5667[68]), .B0(cout_adj_5134), 
          .C0(n87_adj_5565), .D0(d2_adj_5668[68]), .A1(d1_adj_5667[69]), 
          .B1(cout_adj_5134), .C1(n84_adj_5564), .D1(d2_adj_5668[69]), 
          .CIN(n15432), .COUT(n15433), .S0(d2_71__N_490_adj_5684[68]), 
          .S1(d2_71__N_490_adj_5684[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_33 (.A0(d1_adj_5667[66]), .B0(cout_adj_5134), 
          .C0(n93_adj_5567), .D0(d2_adj_5668[66]), .A1(d1_adj_5667[67]), 
          .B1(cout_adj_5134), .C1(n90_adj_5566), .D1(d2_adj_5668[67]), 
          .CIN(n15431), .COUT(n15432), .S0(d2_71__N_490_adj_5684[66]), 
          .S1(d2_71__N_490_adj_5684[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_31 (.A0(d1_adj_5667[64]), .B0(cout_adj_5134), 
          .C0(n99_adj_5569), .D0(d2_adj_5668[64]), .A1(d1_adj_5667[65]), 
          .B1(cout_adj_5134), .C1(n96_adj_5568), .D1(d2_adj_5668[65]), 
          .CIN(n15430), .COUT(n15431), .S0(d2_71__N_490_adj_5684[64]), 
          .S1(d2_71__N_490_adj_5684[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_29 (.A0(d1_adj_5667[62]), .B0(cout_adj_5134), 
          .C0(n105_adj_5571), .D0(d2_adj_5668[62]), .A1(d1_adj_5667[63]), 
          .B1(cout_adj_5134), .C1(n102_adj_5570), .D1(d2_adj_5668[63]), 
          .CIN(n15429), .COUT(n15430), .S0(d2_71__N_490_adj_5684[62]), 
          .S1(d2_71__N_490_adj_5684[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_27 (.A0(d1_adj_5667[60]), .B0(cout_adj_5134), 
          .C0(n111_adj_5573), .D0(d2_adj_5668[60]), .A1(d1_adj_5667[61]), 
          .B1(cout_adj_5134), .C1(n108_adj_5572), .D1(d2_adj_5668[61]), 
          .CIN(n15428), .COUT(n15429), .S0(d2_71__N_490_adj_5684[60]), 
          .S1(d2_71__N_490_adj_5684[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_25 (.A0(d1_adj_5667[58]), .B0(cout_adj_5134), 
          .C0(n117_adj_5575), .D0(d2_adj_5668[58]), .A1(d1_adj_5667[59]), 
          .B1(cout_adj_5134), .C1(n114_adj_5574), .D1(d2_adj_5668[59]), 
          .CIN(n15427), .COUT(n15428), .S0(d2_71__N_490_adj_5684[58]), 
          .S1(d2_71__N_490_adj_5684[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_23 (.A0(d1_adj_5667[56]), .B0(cout_adj_5134), 
          .C0(n123_adj_5577), .D0(d2_adj_5668[56]), .A1(d1_adj_5667[57]), 
          .B1(cout_adj_5134), .C1(n120_adj_5576), .D1(d2_adj_5668[57]), 
          .CIN(n15426), .COUT(n15427), .S0(d2_71__N_490_adj_5684[56]), 
          .S1(d2_71__N_490_adj_5684[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_21 (.A0(d1_adj_5667[54]), .B0(cout_adj_5134), 
          .C0(n129_adj_5579), .D0(d2_adj_5668[54]), .A1(d1_adj_5667[55]), 
          .B1(cout_adj_5134), .C1(n126_adj_5578), .D1(d2_adj_5668[55]), 
          .CIN(n15425), .COUT(n15426), .S0(d2_71__N_490_adj_5684[54]), 
          .S1(d2_71__N_490_adj_5684[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_19 (.A0(d1_adj_5667[52]), .B0(cout_adj_5134), 
          .C0(n135_adj_5581), .D0(d2_adj_5668[52]), .A1(d1_adj_5667[53]), 
          .B1(cout_adj_5134), .C1(n132_adj_5580), .D1(d2_adj_5668[53]), 
          .CIN(n15424), .COUT(n15425), .S0(d2_71__N_490_adj_5684[52]), 
          .S1(d2_71__N_490_adj_5684[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_17 (.A0(d1_adj_5667[50]), .B0(cout_adj_5134), 
          .C0(n141_adj_5583), .D0(d2_adj_5668[50]), .A1(d1_adj_5667[51]), 
          .B1(cout_adj_5134), .C1(n138_adj_5582), .D1(d2_adj_5668[51]), 
          .CIN(n15423), .COUT(n15424), .S0(d2_71__N_490_adj_5684[50]), 
          .S1(d2_71__N_490_adj_5684[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_15 (.A0(d1_adj_5667[48]), .B0(cout_adj_5134), 
          .C0(n147_adj_5585), .D0(d2_adj_5668[48]), .A1(d1_adj_5667[49]), 
          .B1(cout_adj_5134), .C1(n144_adj_5584), .D1(d2_adj_5668[49]), 
          .CIN(n15422), .COUT(n15423), .S0(d2_71__N_490_adj_5684[48]), 
          .S1(d2_71__N_490_adj_5684[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_13 (.A0(d1_adj_5667[46]), .B0(cout_adj_5134), 
          .C0(n153_adj_5587), .D0(d2_adj_5668[46]), .A1(d1_adj_5667[47]), 
          .B1(cout_adj_5134), .C1(n150_adj_5586), .D1(d2_adj_5668[47]), 
          .CIN(n15421), .COUT(n15422), .S0(d2_71__N_490_adj_5684[46]), 
          .S1(d2_71__N_490_adj_5684[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_11 (.A0(d1_adj_5667[44]), .B0(cout_adj_5134), 
          .C0(n159_adj_5589), .D0(d2_adj_5668[44]), .A1(d1_adj_5667[45]), 
          .B1(cout_adj_5134), .C1(n156_adj_5588), .D1(d2_adj_5668[45]), 
          .CIN(n15420), .COUT(n15421), .S0(d2_71__N_490_adj_5684[44]), 
          .S1(d2_71__N_490_adj_5684[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_9 (.A0(d1_adj_5667[42]), .B0(cout_adj_5134), 
          .C0(n165_adj_5591), .D0(d2_adj_5668[42]), .A1(d1_adj_5667[43]), 
          .B1(cout_adj_5134), .C1(n162_adj_5590), .D1(d2_adj_5668[43]), 
          .CIN(n15419), .COUT(n15420), .S0(d2_71__N_490_adj_5684[42]), 
          .S1(d2_71__N_490_adj_5684[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_7 (.A0(d1_adj_5667[40]), .B0(cout_adj_5134), 
          .C0(n171_adj_5593), .D0(d2_adj_5668[40]), .A1(d1_adj_5667[41]), 
          .B1(cout_adj_5134), .C1(n168_adj_5592), .D1(d2_adj_5668[41]), 
          .CIN(n15418), .COUT(n15419), .S0(d2_71__N_490_adj_5684[40]), 
          .S1(d2_71__N_490_adj_5684[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_5 (.A0(d1_adj_5667[38]), .B0(cout_adj_5134), 
          .C0(n177_adj_5595), .D0(d2_adj_5668[38]), .A1(d1_adj_5667[39]), 
          .B1(cout_adj_5134), .C1(n174_adj_5594), .D1(d2_adj_5668[39]), 
          .CIN(n15417), .COUT(n15418), .S0(d2_71__N_490_adj_5684[38]), 
          .S1(d2_71__N_490_adj_5684[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_3 (.A0(d1_adj_5667[36]), .B0(cout_adj_5134), 
          .C0(n183_adj_5597), .D0(d2_adj_5668[36]), .A1(d1_adj_5667[37]), 
          .B1(cout_adj_5134), .C1(n180_adj_5596), .D1(d2_adj_5668[37]), 
          .CIN(n15416), .COUT(n15417), .S0(d2_71__N_490_adj_5684[36]), 
          .S1(d2_71__N_490_adj_5684[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1499_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1499_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1499_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5134), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15416));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1499_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1499_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1499_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1499_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_38 (.A0(d3[71]), .B0(d2[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15412), .S0(n78_adj_5218));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1556_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_36 (.A0(d3[69]), .B0(d2[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[70]), .B1(d2[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15411), .COUT(n15412), .S0(n84_adj_5220), .S1(n81_adj_5219));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_34 (.A0(d3[67]), .B0(d2[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[68]), .B1(d2[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15410), .COUT(n15411), .S0(n90_adj_5222), .S1(n87_adj_5221));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_32 (.A0(d3[65]), .B0(d2[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[66]), .B1(d2[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15409), .COUT(n15410), .S0(n96_adj_5224), .S1(n93_adj_5223));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_30 (.A0(d3[63]), .B0(d2[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[64]), .B1(d2[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15408), .COUT(n15409), .S0(n102_adj_5226), .S1(n99_adj_5225));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_28 (.A0(d3[61]), .B0(d2[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[62]), .B1(d2[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15407), .COUT(n15408), .S0(n108_adj_5228), .S1(n105_adj_5227));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_26 (.A0(d3[59]), .B0(d2[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[60]), .B1(d2[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15406), .COUT(n15407), .S0(n114_adj_5230), .S1(n111_adj_5229));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_24 (.A0(d3[57]), .B0(d2[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[58]), .B1(d2[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15405), .COUT(n15406), .S0(n120_adj_5232), .S1(n117_adj_5231));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_22 (.A0(d3[55]), .B0(d2[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[56]), .B1(d2[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15404), .COUT(n15405), .S0(n126_adj_5234), .S1(n123_adj_5233));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_20 (.A0(d3[53]), .B0(d2[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[54]), .B1(d2[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15403), .COUT(n15404), .S0(n132_adj_5236), .S1(n129_adj_5235));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_18 (.A0(d3[51]), .B0(d2[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[52]), .B1(d2[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15402), .COUT(n15403), .S0(n138_adj_5238), .S1(n135_adj_5237));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_16 (.A0(d3[49]), .B0(d2[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[50]), .B1(d2[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15401), .COUT(n15402), .S0(n144_adj_5240), .S1(n141_adj_5239));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_14 (.A0(d3[47]), .B0(d2[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[48]), .B1(d2[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15400), .COUT(n15401), .S0(n150_adj_5242), .S1(n147_adj_5241));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_12 (.A0(d3[45]), .B0(d2[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[46]), .B1(d2[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15399), .COUT(n15400), .S0(n156_adj_5244), .S1(n153_adj_5243));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_10 (.A0(d3[43]), .B0(d2[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[44]), .B1(d2[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15398), .COUT(n15399), .S0(n162_adj_5246), .S1(n159_adj_5245));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_8 (.A0(d3[41]), .B0(d2[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[42]), .B1(d2[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15397), .COUT(n15398), .S0(n168_adj_5248), .S1(n165_adj_5247));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_6 (.A0(d3[39]), .B0(d2[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[40]), .B1(d2[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15396), .COUT(n15397), .S0(n174_adj_5250), .S1(n171_adj_5249));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_4 (.A0(d3[37]), .B0(d2[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[38]), .B1(d2[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15395), .COUT(n15396), .S0(n180_adj_5252), .S1(n177_adj_5251));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1556_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[36]), .B1(d2[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15395), .S1(n183_adj_5253));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1556_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1556_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1556_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_38 (.A0(d5_adj_5671[71]), .B0(d4_adj_5670[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15394), .S0(n78_adj_2773));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1577_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_36 (.A0(d5_adj_5671[69]), .B0(d4_adj_5670[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[70]), .B1(d4_adj_5670[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15393), .COUT(n15394), .S0(n84_adj_2771), 
          .S1(n81_adj_2772));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_36.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_169 (.A(o_Rx_DV), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[7]), 
         .Z(n17638)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_169.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_163_4_lut (.A(o_Rx_DV), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[7]), 
         .D(o_Rx_Byte[6]), .Z(n17632)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_163_4_lut.init = 16'hf7ff;
    LUT4 i1_2_lut_4_lut (.A(o_Rx_DV), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[7]), 
         .D(o_Rx_Byte[4]), .Z(n16812)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_2_lut_4_lut.init = 16'hf7ff;
    CCU2C _add_1_1577_add_4_34 (.A0(d5_adj_5671[67]), .B0(d4_adj_5670[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[68]), .B1(d4_adj_5670[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15392), .COUT(n15393), .S0(n90_adj_2769), 
          .S1(n87_adj_2770));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_32 (.A0(d5_adj_5671[65]), .B0(d4_adj_5670[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[66]), .B1(d4_adj_5670[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15391), .COUT(n15392), .S0(n96), 
          .S1(n93));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_30 (.A0(d5_adj_5671[63]), .B0(d4_adj_5670[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[64]), .B1(d4_adj_5670[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15390), .COUT(n15391), .S0(n102), 
          .S1(n99));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_28 (.A0(d5_adj_5671[61]), .B0(d4_adj_5670[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[62]), .B1(d4_adj_5670[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15389), .COUT(n15390), .S0(n108), 
          .S1(n105));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_26 (.A0(d5_adj_5671[59]), .B0(d4_adj_5670[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[60]), .B1(d4_adj_5670[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15388), .COUT(n15389), .S0(n114), 
          .S1(n111));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_24 (.A0(d5_adj_5671[57]), .B0(d4_adj_5670[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[58]), .B1(d4_adj_5670[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15387), .COUT(n15388), .S0(n120), 
          .S1(n117));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_22 (.A0(d5_adj_5671[55]), .B0(d4_adj_5670[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[56]), .B1(d4_adj_5670[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15386), .COUT(n15387), .S0(n126), 
          .S1(n123));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_20 (.A0(d5_adj_5671[53]), .B0(d4_adj_5670[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[54]), .B1(d4_adj_5670[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15385), .COUT(n15386), .S0(n132), 
          .S1(n129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_18 (.A0(d5_adj_5671[51]), .B0(d4_adj_5670[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[52]), .B1(d4_adj_5670[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15384), .COUT(n15385), .S0(n138), 
          .S1(n135));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_16 (.A0(d5_adj_5671[49]), .B0(d4_adj_5670[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[50]), .B1(d4_adj_5670[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15383), .COUT(n15384), .S0(n144), 
          .S1(n141));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_14 (.A0(d5_adj_5671[47]), .B0(d4_adj_5670[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[48]), .B1(d4_adj_5670[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15382), .COUT(n15383), .S0(n150), 
          .S1(n147));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_12 (.A0(d5_adj_5671[45]), .B0(d4_adj_5670[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[46]), .B1(d4_adj_5670[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15381), .COUT(n15382), .S0(n156), 
          .S1(n153));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_10 (.A0(d5_adj_5671[43]), .B0(d4_adj_5670[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[44]), .B1(d4_adj_5670[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15380), .COUT(n15381), .S0(n162), 
          .S1(n159));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_8 (.A0(d5_adj_5671[41]), .B0(d4_adj_5670[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[42]), .B1(d4_adj_5670[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15379), .COUT(n15380), .S0(n168_adj_2767), 
          .S1(n165_adj_2768));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_6 (.A0(d5_adj_5671[39]), .B0(d4_adj_5670[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[40]), .B1(d4_adj_5670[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15378), .COUT(n15379), .S0(n174_adj_2765), 
          .S1(n171_adj_2766));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_4 (.A0(d5_adj_5671[37]), .B0(d4_adj_5670[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5671[38]), .B1(d4_adj_5670[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15377), .COUT(n15378), .S0(n180_adj_2763), 
          .S1(n177_adj_2764));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1577_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5_adj_5671[36]), .B1(d4_adj_5670[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15377), .S1(n183));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1577_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1577_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1577_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_37 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n81_adj_5438), .D0(d1_adj_5667[70]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n78_adj_5437), .D1(d1_adj_5667[71]), 
          .CIN(n15375), .S0(d1_71__N_418_adj_5683[70]), .S1(d1_71__N_418_adj_5683[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_35 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n87_adj_5440), .D0(d1_adj_5667[68]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n84_adj_5439), .D1(d1_adj_5667[69]), 
          .CIN(n15374), .COUT(n15375), .S0(d1_71__N_418_adj_5683[68]), 
          .S1(d1_71__N_418_adj_5683[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_33 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n93_adj_5442), .D0(d1_adj_5667[66]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n90_adj_5441), .D1(d1_adj_5667[67]), 
          .CIN(n15373), .COUT(n15374), .S0(d1_71__N_418_adj_5683[66]), 
          .S1(d1_71__N_418_adj_5683[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_31 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n99_adj_5444), .D0(d1_adj_5667[64]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n96_adj_5443), .D1(d1_adj_5667[65]), 
          .CIN(n15372), .COUT(n15373), .S0(d1_71__N_418_adj_5683[64]), 
          .S1(d1_71__N_418_adj_5683[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_29 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n105_adj_5446), .D0(d1_adj_5667[62]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n102_adj_5445), .D1(d1_adj_5667[63]), 
          .CIN(n15371), .COUT(n15372), .S0(d1_71__N_418_adj_5683[62]), 
          .S1(d1_71__N_418_adj_5683[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_27 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n111_adj_5448), .D0(d1_adj_5667[60]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n108_adj_5447), .D1(d1_adj_5667[61]), 
          .CIN(n15370), .COUT(n15371), .S0(d1_71__N_418_adj_5683[60]), 
          .S1(d1_71__N_418_adj_5683[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_25 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n117_adj_5450), .D0(d1_adj_5667[58]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n114_adj_5449), .D1(d1_adj_5667[59]), 
          .CIN(n15369), .COUT(n15370), .S0(d1_71__N_418_adj_5683[58]), 
          .S1(d1_71__N_418_adj_5683[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_23 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n123_adj_5452), .D0(d1_adj_5667[56]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n120_adj_5451), .D1(d1_adj_5667[57]), 
          .CIN(n15368), .COUT(n15369), .S0(d1_71__N_418_adj_5683[56]), 
          .S1(d1_71__N_418_adj_5683[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_21 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n129_adj_5454), .D0(d1_adj_5667[54]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n126_adj_5453), .D1(d1_adj_5667[55]), 
          .CIN(n15367), .COUT(n15368), .S0(d1_71__N_418_adj_5683[54]), 
          .S1(d1_71__N_418_adj_5683[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_19 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n135_adj_5456), .D0(d1_adj_5667[52]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n132_adj_5455), .D1(d1_adj_5667[53]), 
          .CIN(n15366), .COUT(n15367), .S0(d1_71__N_418_adj_5683[52]), 
          .S1(d1_71__N_418_adj_5683[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_17 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n141_adj_5458), .D0(d1_adj_5667[50]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n138_adj_5457), .D1(d1_adj_5667[51]), 
          .CIN(n15365), .COUT(n15366), .S0(d1_71__N_418_adj_5683[50]), 
          .S1(d1_71__N_418_adj_5683[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_15 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n147_adj_5460), .D0(d1_adj_5667[48]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n144_adj_5459), .D1(d1_adj_5667[49]), 
          .CIN(n15364), .COUT(n15365), .S0(d1_71__N_418_adj_5683[48]), 
          .S1(d1_71__N_418_adj_5683[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_13 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n153_adj_5462), .D0(d1_adj_5667[46]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n150_adj_5461), .D1(d1_adj_5667[47]), 
          .CIN(n15363), .COUT(n15364), .S0(d1_71__N_418_adj_5683[46]), 
          .S1(d1_71__N_418_adj_5683[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_11 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n159_adj_5464), .D0(d1_adj_5667[44]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n156_adj_5463), .D1(d1_adj_5667[45]), 
          .CIN(n15362), .COUT(n15363), .S0(d1_71__N_418_adj_5683[44]), 
          .S1(d1_71__N_418_adj_5683[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_9 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n165_adj_5466), .D0(d1_adj_5667[42]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n162_adj_5465), .D1(d1_adj_5667[43]), 
          .CIN(n15361), .COUT(n15362), .S0(d1_71__N_418_adj_5683[42]), 
          .S1(d1_71__N_418_adj_5683[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_7 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n171_adj_5468), .D0(d1_adj_5667[40]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n168_adj_5467), .D1(d1_adj_5667[41]), 
          .CIN(n15360), .COUT(n15361), .S0(d1_71__N_418_adj_5683[40]), 
          .S1(d1_71__N_418_adj_5683[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_5 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n177_adj_5470), .D0(d1_adj_5667[38]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n174_adj_5469), .D1(d1_adj_5667[39]), 
          .CIN(n15359), .COUT(n15360), .S0(d1_71__N_418_adj_5683[38]), 
          .S1(d1_71__N_418_adj_5683[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_3 (.A0(MixerOutCos[11]), .B0(cout_adj_5128), 
          .C0(n183_adj_5472), .D0(d1_adj_5667[36]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5128), .C1(n180_adj_5471), .D1(d1_adj_5667[37]), 
          .CIN(n15358), .COUT(n15359), .S0(d1_71__N_418_adj_5683[36]), 
          .S1(d1_71__N_418_adj_5683[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1502_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1502_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1502_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5128), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15358));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1502_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1502_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1502_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1502_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_37 (.A0(d4[70]), .B0(cout_adj_5127), .C0(n81_adj_5385), 
          .D0(d5[70]), .A1(d4[71]), .B1(cout_adj_5127), .C1(n78_adj_5384), 
          .D1(d5[71]), .CIN(n15353), .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_35 (.A0(d4[68]), .B0(cout_adj_5127), .C0(n87_adj_5387), 
          .D0(d5[68]), .A1(d4[69]), .B1(cout_adj_5127), .C1(n84_adj_5386), 
          .D1(d5[69]), .CIN(n15352), .COUT(n15353), .S0(d5_71__N_706[68]), 
          .S1(d5_71__N_706[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_33 (.A0(d4[66]), .B0(cout_adj_5127), .C0(n93_adj_5389), 
          .D0(d5[66]), .A1(d4[67]), .B1(cout_adj_5127), .C1(n90_adj_5388), 
          .D1(d5[67]), .CIN(n15351), .COUT(n15352), .S0(d5_71__N_706[66]), 
          .S1(d5_71__N_706[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_31 (.A0(d4[64]), .B0(cout_adj_5127), .C0(n99_adj_5391), 
          .D0(d5[64]), .A1(d4[65]), .B1(cout_adj_5127), .C1(n96_adj_5390), 
          .D1(d5[65]), .CIN(n15350), .COUT(n15351), .S0(d5_71__N_706[64]), 
          .S1(d5_71__N_706[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_29 (.A0(d4[62]), .B0(cout_adj_5127), .C0(n105_adj_5393), 
          .D0(d5[62]), .A1(d4[63]), .B1(cout_adj_5127), .C1(n102_adj_5392), 
          .D1(d5[63]), .CIN(n15349), .COUT(n15350), .S0(d5_71__N_706[62]), 
          .S1(d5_71__N_706[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_27 (.A0(d4[60]), .B0(cout_adj_5127), .C0(n111_adj_5395), 
          .D0(d5[60]), .A1(d4[61]), .B1(cout_adj_5127), .C1(n108_adj_5394), 
          .D1(d5[61]), .CIN(n15348), .COUT(n15349), .S0(d5_71__N_706[60]), 
          .S1(d5_71__N_706[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_25 (.A0(d4[58]), .B0(cout_adj_5127), .C0(n117_adj_5397), 
          .D0(d5[58]), .A1(d4[59]), .B1(cout_adj_5127), .C1(n114_adj_5396), 
          .D1(d5[59]), .CIN(n15347), .COUT(n15348), .S0(d5_71__N_706[58]), 
          .S1(d5_71__N_706[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_23 (.A0(d4[56]), .B0(cout_adj_5127), .C0(n123_adj_5399), 
          .D0(d5[56]), .A1(d4[57]), .B1(cout_adj_5127), .C1(n120_adj_5398), 
          .D1(d5[57]), .CIN(n15346), .COUT(n15347), .S0(d5_71__N_706[56]), 
          .S1(d5_71__N_706[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_21 (.A0(d4[54]), .B0(cout_adj_5127), .C0(n129_adj_5401), 
          .D0(d5[54]), .A1(d4[55]), .B1(cout_adj_5127), .C1(n126_adj_5400), 
          .D1(d5[55]), .CIN(n15345), .COUT(n15346), .S0(d5_71__N_706[54]), 
          .S1(d5_71__N_706[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_19 (.A0(d4[52]), .B0(cout_adj_5127), .C0(n135_adj_5403), 
          .D0(d5[52]), .A1(d4[53]), .B1(cout_adj_5127), .C1(n132_adj_5402), 
          .D1(d5[53]), .CIN(n15344), .COUT(n15345), .S0(d5_71__N_706[52]), 
          .S1(d5_71__N_706[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_17 (.A0(d4[50]), .B0(cout_adj_5127), .C0(n141_adj_5405), 
          .D0(d5[50]), .A1(d4[51]), .B1(cout_adj_5127), .C1(n138_adj_5404), 
          .D1(d5[51]), .CIN(n15343), .COUT(n15344), .S0(d5_71__N_706[50]), 
          .S1(d5_71__N_706[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_15 (.A0(d4[48]), .B0(cout_adj_5127), .C0(n147_adj_5407), 
          .D0(d5[48]), .A1(d4[49]), .B1(cout_adj_5127), .C1(n144_adj_5406), 
          .D1(d5[49]), .CIN(n15342), .COUT(n15343), .S0(d5_71__N_706[48]), 
          .S1(d5_71__N_706[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_13 (.A0(d4[46]), .B0(cout_adj_5127), .C0(n153_adj_5409), 
          .D0(d5[46]), .A1(d4[47]), .B1(cout_adj_5127), .C1(n150_adj_5408), 
          .D1(d5[47]), .CIN(n15341), .COUT(n15342), .S0(d5_71__N_706[46]), 
          .S1(d5_71__N_706[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_11 (.A0(d4[44]), .B0(cout_adj_5127), .C0(n159_adj_5411), 
          .D0(d5[44]), .A1(d4[45]), .B1(cout_adj_5127), .C1(n156_adj_5410), 
          .D1(d5[45]), .CIN(n15340), .COUT(n15341), .S0(d5_71__N_706[44]), 
          .S1(d5_71__N_706[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_9 (.A0(d4[42]), .B0(cout_adj_5127), .C0(n165_adj_5413), 
          .D0(d5[42]), .A1(d4[43]), .B1(cout_adj_5127), .C1(n162_adj_5412), 
          .D1(d5[43]), .CIN(n15339), .COUT(n15340), .S0(d5_71__N_706[42]), 
          .S1(d5_71__N_706[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_7 (.A0(d4[40]), .B0(cout_adj_5127), .C0(n171_adj_5415), 
          .D0(d5[40]), .A1(d4[41]), .B1(cout_adj_5127), .C1(n168_adj_5414), 
          .D1(d5[41]), .CIN(n15338), .COUT(n15339), .S0(d5_71__N_706[40]), 
          .S1(d5_71__N_706[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_5 (.A0(d4[38]), .B0(cout_adj_5127), .C0(n177_adj_5417), 
          .D0(d5[38]), .A1(d4[39]), .B1(cout_adj_5127), .C1(n174_adj_5416), 
          .D1(d5[39]), .CIN(n15337), .COUT(n15338), .S0(d5_71__N_706[38]), 
          .S1(d5_71__N_706[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_3 (.A0(d4[36]), .B0(cout_adj_5127), .C0(n183_adj_5419), 
          .D0(d5[36]), .A1(d4[37]), .B1(cout_adj_5127), .C1(n180_adj_5418), 
          .D1(d5[37]), .CIN(n15336), .COUT(n15337), .S0(d5_71__N_706[36]), 
          .S1(d5_71__N_706[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1505_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1505_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1505_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5127), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15336));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1505_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1505_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1505_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1505_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_37 (.A0(d3[70]), .B0(cout_adj_5126), .C0(n81_adj_5343), 
          .D0(d4[70]), .A1(d3[71]), .B1(cout_adj_5126), .C1(n78_adj_5342), 
          .D1(d4[71]), .CIN(n15331), .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_35 (.A0(d3[68]), .B0(cout_adj_5126), .C0(n87_adj_5345), 
          .D0(d4[68]), .A1(d3[69]), .B1(cout_adj_5126), .C1(n84_adj_5344), 
          .D1(d4[69]), .CIN(n15330), .COUT(n15331), .S0(d4_71__N_634[68]), 
          .S1(d4_71__N_634[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_33 (.A0(d3[66]), .B0(cout_adj_5126), .C0(n93_adj_5347), 
          .D0(d4[66]), .A1(d3[67]), .B1(cout_adj_5126), .C1(n90_adj_5346), 
          .D1(d4[67]), .CIN(n15329), .COUT(n15330), .S0(d4_71__N_634[66]), 
          .S1(d4_71__N_634[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_31 (.A0(d3[64]), .B0(cout_adj_5126), .C0(n99_adj_5349), 
          .D0(d4[64]), .A1(d3[65]), .B1(cout_adj_5126), .C1(n96_adj_5348), 
          .D1(d4[65]), .CIN(n15328), .COUT(n15329), .S0(d4_71__N_634[64]), 
          .S1(d4_71__N_634[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_29 (.A0(d3[62]), .B0(cout_adj_5126), .C0(n105_adj_5351), 
          .D0(d4[62]), .A1(d3[63]), .B1(cout_adj_5126), .C1(n102_adj_5350), 
          .D1(d4[63]), .CIN(n15327), .COUT(n15328), .S0(d4_71__N_634[62]), 
          .S1(d4_71__N_634[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_27 (.A0(d3[60]), .B0(cout_adj_5126), .C0(n111_adj_5353), 
          .D0(d4[60]), .A1(d3[61]), .B1(cout_adj_5126), .C1(n108_adj_5352), 
          .D1(d4[61]), .CIN(n15326), .COUT(n15327), .S0(d4_71__N_634[60]), 
          .S1(d4_71__N_634[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_25 (.A0(d3[58]), .B0(cout_adj_5126), .C0(n117_adj_5355), 
          .D0(d4[58]), .A1(d3[59]), .B1(cout_adj_5126), .C1(n114_adj_5354), 
          .D1(d4[59]), .CIN(n15325), .COUT(n15326), .S0(d4_71__N_634[58]), 
          .S1(d4_71__N_634[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_23 (.A0(d3[56]), .B0(cout_adj_5126), .C0(n123_adj_5357), 
          .D0(d4[56]), .A1(d3[57]), .B1(cout_adj_5126), .C1(n120_adj_5356), 
          .D1(d4[57]), .CIN(n15324), .COUT(n15325), .S0(d4_71__N_634[56]), 
          .S1(d4_71__N_634[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_21 (.A0(d3[54]), .B0(cout_adj_5126), .C0(n129_adj_5359), 
          .D0(d4[54]), .A1(d3[55]), .B1(cout_adj_5126), .C1(n126_adj_5358), 
          .D1(d4[55]), .CIN(n15323), .COUT(n15324), .S0(d4_71__N_634[54]), 
          .S1(d4_71__N_634[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_19 (.A0(d3[52]), .B0(cout_adj_5126), .C0(n135_adj_5361), 
          .D0(d4[52]), .A1(d3[53]), .B1(cout_adj_5126), .C1(n132_adj_5360), 
          .D1(d4[53]), .CIN(n15322), .COUT(n15323), .S0(d4_71__N_634[52]), 
          .S1(d4_71__N_634[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_17 (.A0(d3[50]), .B0(cout_adj_5126), .C0(n141_adj_5363), 
          .D0(d4[50]), .A1(d3[51]), .B1(cout_adj_5126), .C1(n138_adj_5362), 
          .D1(d4[51]), .CIN(n15321), .COUT(n15322), .S0(d4_71__N_634[50]), 
          .S1(d4_71__N_634[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_15 (.A0(d3[48]), .B0(cout_adj_5126), .C0(n147_adj_5365), 
          .D0(d4[48]), .A1(d3[49]), .B1(cout_adj_5126), .C1(n144_adj_5364), 
          .D1(d4[49]), .CIN(n15320), .COUT(n15321), .S0(d4_71__N_634[48]), 
          .S1(d4_71__N_634[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_13 (.A0(d3[46]), .B0(cout_adj_5126), .C0(n153_adj_5367), 
          .D0(d4[46]), .A1(d3[47]), .B1(cout_adj_5126), .C1(n150_adj_5366), 
          .D1(d4[47]), .CIN(n15319), .COUT(n15320), .S0(d4_71__N_634[46]), 
          .S1(d4_71__N_634[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_11 (.A0(d3[44]), .B0(cout_adj_5126), .C0(n159_adj_5369), 
          .D0(d4[44]), .A1(d3[45]), .B1(cout_adj_5126), .C1(n156_adj_5368), 
          .D1(d4[45]), .CIN(n15318), .COUT(n15319), .S0(d4_71__N_634[44]), 
          .S1(d4_71__N_634[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_9 (.A0(d3[42]), .B0(cout_adj_5126), .C0(n165_adj_5371), 
          .D0(d4[42]), .A1(d3[43]), .B1(cout_adj_5126), .C1(n162_adj_5370), 
          .D1(d4[43]), .CIN(n15317), .COUT(n15318), .S0(d4_71__N_634[42]), 
          .S1(d4_71__N_634[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_7 (.A0(d3[40]), .B0(cout_adj_5126), .C0(n171_adj_5373), 
          .D0(d4[40]), .A1(d3[41]), .B1(cout_adj_5126), .C1(n168_adj_5372), 
          .D1(d4[41]), .CIN(n15316), .COUT(n15317), .S0(d4_71__N_634[40]), 
          .S1(d4_71__N_634[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_5 (.A0(d3[38]), .B0(cout_adj_5126), .C0(n177_adj_5375), 
          .D0(d4[38]), .A1(d3[39]), .B1(cout_adj_5126), .C1(n174_adj_5374), 
          .D1(d4[39]), .CIN(n15315), .COUT(n15316), .S0(d4_71__N_634[38]), 
          .S1(d4_71__N_634[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_3 (.A0(d3[36]), .B0(cout_adj_5126), .C0(n183_adj_5377), 
          .D0(d4[36]), .A1(d3[37]), .B1(cout_adj_5126), .C1(n180_adj_5376), 
          .D1(d4[37]), .CIN(n15314), .COUT(n15315), .S0(d4_71__N_634[36]), 
          .S1(d4_71__N_634[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1508_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1508_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1508_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5126), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1508_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1508_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1508_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1508_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_37 (.A0(d2[70]), .B0(cout_adj_4837), .C0(n81_adj_5219), 
          .D0(d3[70]), .A1(d2[71]), .B1(cout_adj_4837), .C1(n78_adj_5218), 
          .D1(d3[71]), .CIN(n15309), .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_35 (.A0(d2[68]), .B0(cout_adj_4837), .C0(n87_adj_5221), 
          .D0(d3[68]), .A1(d2[69]), .B1(cout_adj_4837), .C1(n84_adj_5220), 
          .D1(d3[69]), .CIN(n15308), .COUT(n15309), .S0(d3_71__N_562[68]), 
          .S1(d3_71__N_562[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_33 (.A0(d2[66]), .B0(cout_adj_4837), .C0(n93_adj_5223), 
          .D0(d3[66]), .A1(d2[67]), .B1(cout_adj_4837), .C1(n90_adj_5222), 
          .D1(d3[67]), .CIN(n15307), .COUT(n15308), .S0(d3_71__N_562[66]), 
          .S1(d3_71__N_562[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_31 (.A0(d2[64]), .B0(cout_adj_4837), .C0(n99_adj_5225), 
          .D0(d3[64]), .A1(d2[65]), .B1(cout_adj_4837), .C1(n96_adj_5224), 
          .D1(d3[65]), .CIN(n15306), .COUT(n15307), .S0(d3_71__N_562[64]), 
          .S1(d3_71__N_562[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_29 (.A0(d2[62]), .B0(cout_adj_4837), .C0(n105_adj_5227), 
          .D0(d3[62]), .A1(d2[63]), .B1(cout_adj_4837), .C1(n102_adj_5226), 
          .D1(d3[63]), .CIN(n15305), .COUT(n15306), .S0(d3_71__N_562[62]), 
          .S1(d3_71__N_562[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_27 (.A0(d2[60]), .B0(cout_adj_4837), .C0(n111_adj_5229), 
          .D0(d3[60]), .A1(d2[61]), .B1(cout_adj_4837), .C1(n108_adj_5228), 
          .D1(d3[61]), .CIN(n15304), .COUT(n15305), .S0(d3_71__N_562[60]), 
          .S1(d3_71__N_562[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_25 (.A0(d2[58]), .B0(cout_adj_4837), .C0(n117_adj_5231), 
          .D0(d3[58]), .A1(d2[59]), .B1(cout_adj_4837), .C1(n114_adj_5230), 
          .D1(d3[59]), .CIN(n15303), .COUT(n15304), .S0(d3_71__N_562[58]), 
          .S1(d3_71__N_562[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_23 (.A0(d2[56]), .B0(cout_adj_4837), .C0(n123_adj_5233), 
          .D0(d3[56]), .A1(d2[57]), .B1(cout_adj_4837), .C1(n120_adj_5232), 
          .D1(d3[57]), .CIN(n15302), .COUT(n15303), .S0(d3_71__N_562[56]), 
          .S1(d3_71__N_562[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_21 (.A0(d2[54]), .B0(cout_adj_4837), .C0(n129_adj_5235), 
          .D0(d3[54]), .A1(d2[55]), .B1(cout_adj_4837), .C1(n126_adj_5234), 
          .D1(d3[55]), .CIN(n15301), .COUT(n15302), .S0(d3_71__N_562[54]), 
          .S1(d3_71__N_562[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_19 (.A0(d2[52]), .B0(cout_adj_4837), .C0(n135_adj_5237), 
          .D0(d3[52]), .A1(d2[53]), .B1(cout_adj_4837), .C1(n132_adj_5236), 
          .D1(d3[53]), .CIN(n15300), .COUT(n15301), .S0(d3_71__N_562[52]), 
          .S1(d3_71__N_562[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_17 (.A0(d2[50]), .B0(cout_adj_4837), .C0(n141_adj_5239), 
          .D0(d3[50]), .A1(d2[51]), .B1(cout_adj_4837), .C1(n138_adj_5238), 
          .D1(d3[51]), .CIN(n15299), .COUT(n15300), .S0(d3_71__N_562[50]), 
          .S1(d3_71__N_562[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_15 (.A0(d2[48]), .B0(cout_adj_4837), .C0(n147_adj_5241), 
          .D0(d3[48]), .A1(d2[49]), .B1(cout_adj_4837), .C1(n144_adj_5240), 
          .D1(d3[49]), .CIN(n15298), .COUT(n15299), .S0(d3_71__N_562[48]), 
          .S1(d3_71__N_562[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_13 (.A0(d2[46]), .B0(cout_adj_4837), .C0(n153_adj_5243), 
          .D0(d3[46]), .A1(d2[47]), .B1(cout_adj_4837), .C1(n150_adj_5242), 
          .D1(d3[47]), .CIN(n15297), .COUT(n15298), .S0(d3_71__N_562[46]), 
          .S1(d3_71__N_562[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_11 (.A0(d2[44]), .B0(cout_adj_4837), .C0(n159_adj_5245), 
          .D0(d3[44]), .A1(d2[45]), .B1(cout_adj_4837), .C1(n156_adj_5244), 
          .D1(d3[45]), .CIN(n15296), .COUT(n15297), .S0(d3_71__N_562[44]), 
          .S1(d3_71__N_562[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_9 (.A0(d2[42]), .B0(cout_adj_4837), .C0(n165_adj_5247), 
          .D0(d3[42]), .A1(d2[43]), .B1(cout_adj_4837), .C1(n162_adj_5246), 
          .D1(d3[43]), .CIN(n15295), .COUT(n15296), .S0(d3_71__N_562[42]), 
          .S1(d3_71__N_562[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_7 (.A0(d2[40]), .B0(cout_adj_4837), .C0(n171_adj_5249), 
          .D0(d3[40]), .A1(d2[41]), .B1(cout_adj_4837), .C1(n168_adj_5248), 
          .D1(d3[41]), .CIN(n15294), .COUT(n15295), .S0(d3_71__N_562[40]), 
          .S1(d3_71__N_562[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_5 (.A0(d2[38]), .B0(cout_adj_4837), .C0(n177_adj_5251), 
          .D0(d3[38]), .A1(d2[39]), .B1(cout_adj_4837), .C1(n174_adj_5250), 
          .D1(d3[39]), .CIN(n15293), .COUT(n15294), .S0(d3_71__N_562[38]), 
          .S1(d3_71__N_562[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_3 (.A0(d2[36]), .B0(cout_adj_4837), .C0(n183_adj_5253), 
          .D0(d3[36]), .A1(d2[37]), .B1(cout_adj_4837), .C1(n180_adj_5252), 
          .D1(d3[37]), .CIN(n15292), .COUT(n15293), .S0(d3_71__N_562[36]), 
          .S1(d3_71__N_562[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1511_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1511_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1511_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4837), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15292));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1511_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1511_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1511_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1511_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_38 (.A0(d1_adj_5667[71]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15288), .S0(n78_adj_5437));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1565_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_36 (.A0(d1_adj_5667[69]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[70]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15287), .COUT(n15288), .S0(n84_adj_5439), 
          .S1(n81_adj_5438));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_34 (.A0(d1_adj_5667[67]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[68]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15286), .COUT(n15287), .S0(n90_adj_5441), 
          .S1(n87_adj_5440));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_32 (.A0(d1_adj_5667[65]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[66]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15285), .COUT(n15286), .S0(n96_adj_5443), 
          .S1(n93_adj_5442));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_22 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15745), .COUT(n15746));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_20 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15744), .COUT(n15745));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_18 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15743), .COUT(n15744));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_16 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15742), .COUT(n15743));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_14 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15741), .COUT(n15742));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_12 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15740), .COUT(n15741));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_10 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15739), .COUT(n15740));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_8 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15738), .COUT(n15739));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_6 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15737), .COUT(n15738));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_4 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15736), .COUT(n15737));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15736));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1583_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1583_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_38 (.A0(d_d_tmp_adj_5666[71]), .B0(d_tmp_adj_5665[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15735), .S0(n78_adj_5052));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1586_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_36 (.A0(d_d_tmp_adj_5666[69]), .B0(d_tmp_adj_5665[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[70]), .B1(d_tmp_adj_5665[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15734), .COUT(n15735), .S0(n84_adj_5054), 
          .S1(n81_adj_5053));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_34 (.A0(d_d_tmp_adj_5666[67]), .B0(d_tmp_adj_5665[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[68]), .B1(d_tmp_adj_5665[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15733), .COUT(n15734), .S0(n90_adj_5056), 
          .S1(n87_adj_5055));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_32 (.A0(d_d_tmp_adj_5666[65]), .B0(d_tmp_adj_5665[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[66]), .B1(d_tmp_adj_5665[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15732), .COUT(n15733), .S0(n96_adj_5058), 
          .S1(n93_adj_5057));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_30 (.A0(d_d_tmp_adj_5666[63]), .B0(d_tmp_adj_5665[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[64]), .B1(d_tmp_adj_5665[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15731), .COUT(n15732), .S0(n102_adj_5060), 
          .S1(n99_adj_5059));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_28 (.A0(d_d_tmp_adj_5666[61]), .B0(d_tmp_adj_5665[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[62]), .B1(d_tmp_adj_5665[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15730), .COUT(n15731), .S0(n108_adj_5062), 
          .S1(n105_adj_5061));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_26 (.A0(d_d_tmp_adj_5666[59]), .B0(d_tmp_adj_5665[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[60]), .B1(d_tmp_adj_5665[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15729), .COUT(n15730), .S0(n114_adj_5064), 
          .S1(n111_adj_5063));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_24 (.A0(d_d_tmp_adj_5666[57]), .B0(d_tmp_adj_5665[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[58]), .B1(d_tmp_adj_5665[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15728), .COUT(n15729), .S0(n120_adj_5066), 
          .S1(n117_adj_5065));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_22 (.A0(d_d_tmp_adj_5666[55]), .B0(d_tmp_adj_5665[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[56]), .B1(d_tmp_adj_5665[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15727), .COUT(n15728), .S0(n126_adj_5068), 
          .S1(n123_adj_5067));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_20 (.A0(d_d_tmp_adj_5666[53]), .B0(d_tmp_adj_5665[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[54]), .B1(d_tmp_adj_5665[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15726), .COUT(n15727), .S0(n132_adj_5070), 
          .S1(n129_adj_5069));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_18 (.A0(d_d_tmp_adj_5666[51]), .B0(d_tmp_adj_5665[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[52]), .B1(d_tmp_adj_5665[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15725), .COUT(n15726), .S0(n138_adj_5072), 
          .S1(n135_adj_5071));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_16 (.A0(d_d_tmp_adj_5666[49]), .B0(d_tmp_adj_5665[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[50]), .B1(d_tmp_adj_5665[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15724), .COUT(n15725), .S0(n144_adj_5074), 
          .S1(n141_adj_5073));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_14 (.A0(d_d_tmp_adj_5666[47]), .B0(d_tmp_adj_5665[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[48]), .B1(d_tmp_adj_5665[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15723), .COUT(n15724), .S0(n150_adj_5076), 
          .S1(n147_adj_5075));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_12 (.A0(d_d_tmp_adj_5666[45]), .B0(d_tmp_adj_5665[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[46]), .B1(d_tmp_adj_5665[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15722), .COUT(n15723), .S0(n156_adj_5078), 
          .S1(n153_adj_5077));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_10 (.A0(d_d_tmp_adj_5666[43]), .B0(d_tmp_adj_5665[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[44]), .B1(d_tmp_adj_5665[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15721), .COUT(n15722), .S0(n162_adj_5080), 
          .S1(n159_adj_5079));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_8 (.A0(d_d_tmp_adj_5666[41]), .B0(d_tmp_adj_5665[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[42]), .B1(d_tmp_adj_5665[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15720), .COUT(n15721), .S0(n168_adj_5082), 
          .S1(n165_adj_5081));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_6 (.A0(d_d_tmp_adj_5666[39]), .B0(d_tmp_adj_5665[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[40]), .B1(d_tmp_adj_5665[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15719), .COUT(n15720), .S0(n174_adj_5084), 
          .S1(n171_adj_5083));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_4 (.A0(d_d_tmp_adj_5666[37]), .B0(d_tmp_adj_5665[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5666[38]), .B1(d_tmp_adj_5665[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15718), .COUT(n15719), .S0(n180_adj_5086), 
          .S1(n177_adj_5085));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5666[36]), .B1(d_tmp_adj_5665[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15718), .S1(n183_adj_5087));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1586_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1586_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_20 (.A0(n912), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15717), .S0(d_out_d_11__N_2335[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_20.INIT0 = 16'h555f;
    defparam _add_1_1589_add_4_20.INIT1 = 16'h0000;
    defparam _add_1_1589_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_18 (.A0(ISquare[31]), .B0(n914), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n913), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15716), .COUT(n15717));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_16 (.A0(n916), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n915), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15715), .COUT(n15716));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1589_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_14 (.A0(d_out_d_11__N_1874[17]), .B0(n918), 
          .C0(GND_net), .D0(VCC_net), .A1(ISquare[31]), .B1(n17642), 
          .C1(n917), .D1(VCC_net), .CIN(n15714), .COUT(n15715));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_1589_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_12 (.A0(d_out_d_11__N_1878[17]), .B0(n920), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n919), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15713), .COUT(n15714));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_10 (.A0(d_out_d_11__N_1882[17]), .B0(n922), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n921), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15712), .COUT(n15713));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_8 (.A0(d_out_d_11__N_1886[17]), .B0(n924), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n923), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15711), .COUT(n15712));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_6 (.A0(d_out_d_11__N_1890[17]), .B0(n926), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n925), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15710), .COUT(n15711));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1589_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_4 (.A0(d_out_d_11__N_1892[17]), .B0(ISquare[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1892[17]), .B1(n927), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15709), .COUT(n15710));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1589_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15709));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[15:27])
    defparam _add_1_1589_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1589_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1589_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_38 (.A0(d_d7[35]), .B0(d7[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15708), .S0(d8_71__N_1603[35]), .S1(cout_adj_5088));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1592_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_36 (.A0(d_d7[33]), .B0(d7[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[34]), .B1(d7[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15707), .COUT(n15708), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_34 (.A0(d_d7[31]), .B0(d7[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[32]), .B1(d7[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15706), .COUT(n15707), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_32 (.A0(d_d7[29]), .B0(d7[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[30]), .B1(d7[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15705), .COUT(n15706), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_30 (.A0(d_d7[27]), .B0(d7[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[28]), .B1(d7[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15704), .COUT(n15705), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_28 (.A0(d_d7[25]), .B0(d7[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[26]), .B1(d7[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15703), .COUT(n15704), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_26 (.A0(d_d7[23]), .B0(d7[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[24]), .B1(d7[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15702), .COUT(n15703), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_24 (.A0(d_d7[21]), .B0(d7[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[22]), .B1(d7[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15701), .COUT(n15702), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_22 (.A0(d_d7[19]), .B0(d7[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[20]), .B1(d7[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15700), .COUT(n15701), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_20 (.A0(d_d7[17]), .B0(d7[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[18]), .B1(d7[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15699), .COUT(n15700), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_18 (.A0(d_d7[15]), .B0(d7[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[16]), .B1(d7[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15698), .COUT(n15699), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_16 (.A0(d_d7[13]), .B0(d7[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[14]), .B1(d7[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15697), .COUT(n15698), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_14 (.A0(d_d7[11]), .B0(d7[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[12]), .B1(d7[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15696), .COUT(n15697), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_12 (.A0(d_d7[9]), .B0(d7[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[10]), .B1(d7[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15695), .COUT(n15696), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_10 (.A0(d_d7[7]), .B0(d7[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[8]), .B1(d7[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15694), .COUT(n15695), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_8 (.A0(d_d7[5]), .B0(d7[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[6]), .B1(d7[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15693), .COUT(n15694), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_6 (.A0(d_d7[3]), .B0(d7[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[4]), .B1(d7[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15692), .COUT(n15693), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_4 (.A0(d_d7[1]), .B0(d7[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[2]), .B1(d7[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15691), .COUT(n15692), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[0]), .B1(d7[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15691), .S1(d8_71__N_1603[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1592_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1592_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_38 (.A0(d_d6[71]), .B0(d6[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15690), .S0(n78_adj_4925));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1640_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_36 (.A0(d_d6[69]), .B0(d6[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[70]), .B1(d6[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15689), .COUT(n15690), .S0(n84_adj_4927), .S1(n81_adj_4926));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_34 (.A0(d_d6[67]), .B0(d6[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[68]), .B1(d6[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15688), .COUT(n15689), .S0(n90_adj_4929), .S1(n87_adj_4928));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_32 (.A0(d_d6[65]), .B0(d6[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[66]), .B1(d6[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15687), .COUT(n15688), .S0(n96_adj_4931), .S1(n93_adj_4930));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_30 (.A0(d_d6[63]), .B0(d6[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[64]), .B1(d6[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15686), .COUT(n15687), .S0(n102_adj_4933), .S1(n99_adj_4932));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_28 (.A0(d_d6[61]), .B0(d6[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[62]), .B1(d6[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15685), .COUT(n15686), .S0(n108_adj_4935), .S1(n105_adj_4934));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_26 (.A0(d_d6[59]), .B0(d6[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[60]), .B1(d6[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15684), .COUT(n15685), .S0(n114_adj_4937), .S1(n111_adj_4936));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_24 (.A0(d_d6[57]), .B0(d6[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[58]), .B1(d6[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15683), .COUT(n15684), .S0(n120_adj_4939), .S1(n117_adj_4938));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_22 (.A0(d_d6[55]), .B0(d6[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[56]), .B1(d6[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15682), .COUT(n15683), .S0(n126_adj_4941), .S1(n123_adj_4940));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_20 (.A0(d_d6[53]), .B0(d6[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[54]), .B1(d6[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15681), .COUT(n15682), .S0(n132_adj_4943), .S1(n129_adj_4942));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_18 (.A0(d_d6[51]), .B0(d6[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[52]), .B1(d6[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15680), .COUT(n15681), .S0(n138_adj_4945), .S1(n135_adj_4944));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_16 (.A0(d_d6[49]), .B0(d6[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[50]), .B1(d6[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15679), .COUT(n15680), .S0(n144_adj_4947), .S1(n141_adj_4946));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_16.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i1 (.D(n318), .CK(clk_80mhz), .Q(phase_accum_adj_5658[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_1640_add_4_14 (.A0(d_d6[47]), .B0(d6[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[48]), .B1(d6[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15678), .COUT(n15679), .S0(n150_adj_4949), .S1(n147_adj_4948));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_12 (.A0(d_d6[45]), .B0(d6[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[46]), .B1(d6[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15677), .COUT(n15678), .S0(n156_adj_4951), .S1(n153_adj_4950));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_10 (.A0(d_d6[43]), .B0(d6[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[44]), .B1(d6[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15676), .COUT(n15677), .S0(n162_adj_4953), .S1(n159_adj_4952));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_8 (.A0(d_d6[41]), .B0(d6[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[42]), .B1(d6[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15675), .COUT(n15676), .S0(n168_adj_4955), .S1(n165_adj_4954));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_6 (.A0(d_d6[39]), .B0(d6[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[40]), .B1(d6[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15674), .COUT(n15675), .S0(n174_adj_4957), .S1(n171_adj_4956));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_4 (.A0(d_d6[37]), .B0(d6[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[38]), .B1(d6[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15673), .COUT(n15674), .S0(n180_adj_4959), .S1(n177_adj_4958));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1640_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1640_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[36]), .B1(d6[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15673), .S1(n183_adj_4960));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1640_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1640_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1640_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1640_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_38 (.A0(d_d_tmp[71]), .B0(d_tmp[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15672), .S0(n78_adj_4961));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1643_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_36 (.A0(d_d_tmp[69]), .B0(d_tmp[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[70]), .B1(d_tmp[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15671), .COUT(n15672), .S0(n84_adj_4963), 
          .S1(n81_adj_4962));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_34 (.A0(d_d_tmp[67]), .B0(d_tmp[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[68]), .B1(d_tmp[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15670), .COUT(n15671), .S0(n90_adj_4965), 
          .S1(n87_adj_4964));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_32 (.A0(d_d_tmp[65]), .B0(d_tmp[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[66]), .B1(d_tmp[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15669), .COUT(n15670), .S0(n96_adj_4967), 
          .S1(n93_adj_4966));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_30 (.A0(d_d_tmp[63]), .B0(d_tmp[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[64]), .B1(d_tmp[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15668), .COUT(n15669), .S0(n102_adj_4969), 
          .S1(n99_adj_4968));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_28 (.A0(d_d_tmp[61]), .B0(d_tmp[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[62]), .B1(d_tmp[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15667), .COUT(n15668), .S0(n108_adj_4971), 
          .S1(n105_adj_4970));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_26 (.A0(d_d_tmp[59]), .B0(d_tmp[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[60]), .B1(d_tmp[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15666), .COUT(n15667), .S0(n114_adj_4973), 
          .S1(n111_adj_4972));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_24 (.A0(d_d_tmp[57]), .B0(d_tmp[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[58]), .B1(d_tmp[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15665), .COUT(n15666), .S0(n120_adj_4975), 
          .S1(n117_adj_4974));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_22 (.A0(d_d_tmp[55]), .B0(d_tmp[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[56]), .B1(d_tmp[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15664), .COUT(n15665), .S0(n126_adj_4977), 
          .S1(n123_adj_4976));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_20 (.A0(d_d_tmp[53]), .B0(d_tmp[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[54]), .B1(d_tmp[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15663), .COUT(n15664), .S0(n132_adj_4979), 
          .S1(n129_adj_4978));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_18 (.A0(d_d_tmp[51]), .B0(d_tmp[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[52]), .B1(d_tmp[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15662), .COUT(n15663), .S0(n138_adj_4981), 
          .S1(n135_adj_4980));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_16 (.A0(d_d_tmp[49]), .B0(d_tmp[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[50]), .B1(d_tmp[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15661), .COUT(n15662), .S0(n144_adj_4983), 
          .S1(n141_adj_4982));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_14 (.A0(d_d_tmp[47]), .B0(d_tmp[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[48]), .B1(d_tmp[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15660), .COUT(n15661), .S0(n150_adj_4985), 
          .S1(n147_adj_4984));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_12 (.A0(d_d_tmp[45]), .B0(d_tmp[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[46]), .B1(d_tmp[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15659), .COUT(n15660), .S0(n156_adj_4987), 
          .S1(n153_adj_4986));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_10 (.A0(d_d_tmp[43]), .B0(d_tmp[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[44]), .B1(d_tmp[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15658), .COUT(n15659), .S0(n162_adj_4989), 
          .S1(n159_adj_4988));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_8 (.A0(d_d_tmp[41]), .B0(d_tmp[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[42]), .B1(d_tmp[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15657), .COUT(n15658), .S0(n168_adj_4991), 
          .S1(n165_adj_4990));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_6 (.A0(d_d_tmp[39]), .B0(d_tmp[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[40]), .B1(d_tmp[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15656), .COUT(n15657), .S0(n174_adj_4993), 
          .S1(n171_adj_4992));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_4 (.A0(d_d_tmp[37]), .B0(d_tmp[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[38]), .B1(d_tmp[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15655), .COUT(n15656), .S0(n180_adj_4995), 
          .S1(n177_adj_4994));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1643_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1643_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[36]), .B1(d_tmp[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15655), .S1(n183_adj_4996));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1643_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1643_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1643_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1643_add_4_2.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_64 (.A0(phase_inc_carrGen1[62]), .B0(phase_accum[62]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[63]), .B1(phase_accum[63]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15653), .S0(n135_adj_4537), 
          .S1(n132_adj_4538));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_64.INIT0 = 16'h666a;
    defparam phase_accum_add_4_64.INIT1 = 16'h666a;
    defparam phase_accum_add_4_64.INJECT1_0 = "NO";
    defparam phase_accum_add_4_64.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_62 (.A0(phase_inc_carrGen1[60]), .B0(phase_accum[60]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[61]), .B1(phase_accum[61]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15652), .COUT(n15653), .S0(n141_adj_4535), 
          .S1(n138_adj_4536));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_62.INIT0 = 16'h666a;
    defparam phase_accum_add_4_62.INIT1 = 16'h666a;
    defparam phase_accum_add_4_62.INJECT1_0 = "NO";
    defparam phase_accum_add_4_62.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_60 (.A0(phase_inc_carrGen1[58]), .B0(phase_accum[58]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[59]), .B1(phase_accum[59]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15651), .COUT(n15652), .S0(n147_adj_4533), 
          .S1(n144_adj_4534));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_60.INIT0 = 16'h666a;
    defparam phase_accum_add_4_60.INIT1 = 16'h666a;
    defparam phase_accum_add_4_60.INJECT1_0 = "NO";
    defparam phase_accum_add_4_60.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_58 (.A0(phase_inc_carrGen1[56]), .B0(phase_accum[56]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[57]), .B1(phase_accum[57]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15650), .COUT(n15651), .S0(n153_adj_4531), 
          .S1(n150_adj_4532));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_58.INIT0 = 16'h666a;
    defparam phase_accum_add_4_58.INIT1 = 16'h666a;
    defparam phase_accum_add_4_58.INJECT1_0 = "NO";
    defparam phase_accum_add_4_58.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_56 (.A0(phase_inc_carrGen1[54]), .B0(phase_accum_adj_5658[54]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[55]), .B1(phase_accum_adj_5658[55]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15649), .COUT(n15650), .S0(n159_adj_4529), 
          .S1(n156_adj_4530));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_56.INIT0 = 16'h666a;
    defparam phase_accum_add_4_56.INIT1 = 16'h666a;
    defparam phase_accum_add_4_56.INJECT1_0 = "NO";
    defparam phase_accum_add_4_56.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_54 (.A0(phase_inc_carrGen1[52]), .B0(phase_accum_adj_5658[52]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[53]), .B1(phase_accum_adj_5658[53]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15648), .COUT(n15649), .S0(n165_adj_4527), 
          .S1(n162_adj_4528));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_54.INIT0 = 16'h666a;
    defparam phase_accum_add_4_54.INIT1 = 16'h666a;
    defparam phase_accum_add_4_54.INJECT1_0 = "NO";
    defparam phase_accum_add_4_54.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_52 (.A0(phase_inc_carrGen1[50]), .B0(phase_accum_adj_5658[50]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[51]), .B1(phase_accum_adj_5658[51]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15647), .COUT(n15648), .S0(n171_adj_4525), 
          .S1(n168_adj_4526));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_52.INIT0 = 16'h666a;
    defparam phase_accum_add_4_52.INIT1 = 16'h666a;
    defparam phase_accum_add_4_52.INJECT1_0 = "NO";
    defparam phase_accum_add_4_52.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_50 (.A0(phase_inc_carrGen1[48]), .B0(phase_accum_adj_5658[48]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[49]), .B1(phase_accum_adj_5658[49]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15646), .COUT(n15647), .S0(n177_adj_4523), 
          .S1(n174_adj_4524));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_50.INIT0 = 16'h666a;
    defparam phase_accum_add_4_50.INIT1 = 16'h666a;
    defparam phase_accum_add_4_50.INJECT1_0 = "NO";
    defparam phase_accum_add_4_50.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_48 (.A0(phase_inc_carrGen1[46]), .B0(phase_accum_adj_5658[46]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[47]), .B1(phase_accum_adj_5658[47]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15645), .COUT(n15646), .S0(n183_adj_4521), 
          .S1(n180_adj_4522));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_48.INIT0 = 16'h666a;
    defparam phase_accum_add_4_48.INIT1 = 16'h666a;
    defparam phase_accum_add_4_48.INJECT1_0 = "NO";
    defparam phase_accum_add_4_48.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_46 (.A0(phase_inc_carrGen1[44]), .B0(phase_accum_adj_5658[44]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[45]), .B1(phase_accum_adj_5658[45]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15644), .COUT(n15645), .S0(n189), 
          .S1(n186));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_46.INIT0 = 16'h666a;
    defparam phase_accum_add_4_46.INIT1 = 16'h666a;
    defparam phase_accum_add_4_46.INJECT1_0 = "NO";
    defparam phase_accum_add_4_46.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_44 (.A0(phase_inc_carrGen1[42]), .B0(phase_accum_adj_5658[42]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[43]), .B1(phase_accum_adj_5658[43]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15643), .COUT(n15644), .S0(n195), 
          .S1(n192));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_44.INIT0 = 16'h666a;
    defparam phase_accum_add_4_44.INIT1 = 16'h666a;
    defparam phase_accum_add_4_44.INJECT1_0 = "NO";
    defparam phase_accum_add_4_44.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_42 (.A0(phase_inc_carrGen1[40]), .B0(phase_accum_adj_5658[40]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[41]), .B1(phase_accum_adj_5658[41]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15642), .COUT(n15643), .S0(n201), 
          .S1(n198));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_42.INIT0 = 16'h666a;
    defparam phase_accum_add_4_42.INIT1 = 16'h666a;
    defparam phase_accum_add_4_42.INJECT1_0 = "NO";
    defparam phase_accum_add_4_42.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_40 (.A0(phase_inc_carrGen1[38]), .B0(phase_accum_adj_5658[38]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[39]), .B1(phase_accum_adj_5658[39]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15641), .COUT(n15642), .S0(n207), 
          .S1(n204));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_40.INIT0 = 16'h666a;
    defparam phase_accum_add_4_40.INIT1 = 16'h666a;
    defparam phase_accum_add_4_40.INJECT1_0 = "NO";
    defparam phase_accum_add_4_40.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_38 (.A0(phase_inc_carrGen1[36]), .B0(phase_accum_adj_5658[36]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[37]), .B1(phase_accum_adj_5658[37]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15640), .COUT(n15641), .S0(n213), 
          .S1(n210));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_38.INIT0 = 16'h666a;
    defparam phase_accum_add_4_38.INIT1 = 16'h666a;
    defparam phase_accum_add_4_38.INJECT1_0 = "NO";
    defparam phase_accum_add_4_38.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_36 (.A0(phase_inc_carrGen1[34]), .B0(phase_accum_adj_5658[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[35]), .B1(phase_accum_adj_5658[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15639), .COUT(n15640), .S0(n219), 
          .S1(n216));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_36.INIT0 = 16'h666a;
    defparam phase_accum_add_4_36.INIT1 = 16'h666a;
    defparam phase_accum_add_4_36.INJECT1_0 = "NO";
    defparam phase_accum_add_4_36.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_34 (.A0(phase_inc_carrGen1[32]), .B0(phase_accum_adj_5658[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[33]), .B1(phase_accum_adj_5658[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15638), .COUT(n15639), .S0(n225), 
          .S1(n222));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_34.INIT0 = 16'h666a;
    defparam phase_accum_add_4_34.INIT1 = 16'h666a;
    defparam phase_accum_add_4_34.INJECT1_0 = "NO";
    defparam phase_accum_add_4_34.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_32 (.A0(phase_inc_carrGen1[30]), .B0(phase_accum_adj_5658[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[31]), .B1(phase_accum_adj_5658[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15637), .COUT(n15638), .S0(n231), 
          .S1(n228));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_32.INIT0 = 16'h666a;
    defparam phase_accum_add_4_32.INIT1 = 16'h666a;
    defparam phase_accum_add_4_32.INJECT1_0 = "NO";
    defparam phase_accum_add_4_32.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_30 (.A0(phase_inc_carrGen1[28]), .B0(phase_accum_adj_5658[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[29]), .B1(phase_accum_adj_5658[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15636), .COUT(n15637), .S0(n237), 
          .S1(n234));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_30.INIT0 = 16'h666a;
    defparam phase_accum_add_4_30.INIT1 = 16'h666a;
    defparam phase_accum_add_4_30.INJECT1_0 = "NO";
    defparam phase_accum_add_4_30.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_28 (.A0(phase_inc_carrGen1[26]), .B0(phase_accum_adj_5658[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[27]), .B1(phase_accum_adj_5658[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15635), .COUT(n15636), .S0(n243), 
          .S1(n240));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_28.INIT0 = 16'h666a;
    defparam phase_accum_add_4_28.INIT1 = 16'h666a;
    defparam phase_accum_add_4_28.INJECT1_0 = "NO";
    defparam phase_accum_add_4_28.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_26 (.A0(phase_inc_carrGen1[24]), .B0(phase_accum_adj_5658[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[25]), .B1(phase_accum_adj_5658[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15634), .COUT(n15635), .S0(n249), 
          .S1(n246));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_26.INIT0 = 16'h666a;
    defparam phase_accum_add_4_26.INIT1 = 16'h666a;
    defparam phase_accum_add_4_26.INJECT1_0 = "NO";
    defparam phase_accum_add_4_26.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_24 (.A0(phase_inc_carrGen1[22]), .B0(phase_accum_adj_5658[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[23]), .B1(phase_accum_adj_5658[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15633), .COUT(n15634), .S0(n255), 
          .S1(n252));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_24.INIT0 = 16'h666a;
    defparam phase_accum_add_4_24.INIT1 = 16'h666a;
    defparam phase_accum_add_4_24.INJECT1_0 = "NO";
    defparam phase_accum_add_4_24.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_22 (.A0(phase_inc_carrGen1[20]), .B0(phase_accum_adj_5658[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[21]), .B1(phase_accum_adj_5658[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15632), .COUT(n15633), .S0(n261), 
          .S1(n258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_22.INIT0 = 16'h666a;
    defparam phase_accum_add_4_22.INIT1 = 16'h666a;
    defparam phase_accum_add_4_22.INJECT1_0 = "NO";
    defparam phase_accum_add_4_22.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_20 (.A0(phase_inc_carrGen1[18]), .B0(phase_accum_adj_5658[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[19]), .B1(phase_accum_adj_5658[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15631), .COUT(n15632), .S0(n267), 
          .S1(n264));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_20.INIT0 = 16'h666a;
    defparam phase_accum_add_4_20.INIT1 = 16'h666a;
    defparam phase_accum_add_4_20.INJECT1_0 = "NO";
    defparam phase_accum_add_4_20.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_18 (.A0(phase_inc_carrGen1[16]), .B0(phase_accum_adj_5658[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[17]), .B1(phase_accum_adj_5658[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15630), .COUT(n15631), .S0(n273), 
          .S1(n270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_18.INIT0 = 16'h666a;
    defparam phase_accum_add_4_18.INIT1 = 16'h666a;
    defparam phase_accum_add_4_18.INJECT1_0 = "NO";
    defparam phase_accum_add_4_18.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_16 (.A0(phase_inc_carrGen1[14]), .B0(phase_accum_adj_5658[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[15]), .B1(phase_accum_adj_5658[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15629), .COUT(n15630), .S0(n279), 
          .S1(n276));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_16.INIT0 = 16'h666a;
    defparam phase_accum_add_4_16.INIT1 = 16'h666a;
    defparam phase_accum_add_4_16.INJECT1_0 = "NO";
    defparam phase_accum_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_14 (.A0(phase_inc_carrGen1[12]), .B0(phase_accum_adj_5658[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[13]), .B1(phase_accum_adj_5658[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15628), .COUT(n15629), .S0(n285), 
          .S1(n282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_14.INIT0 = 16'h666a;
    defparam phase_accum_add_4_14.INIT1 = 16'h666a;
    defparam phase_accum_add_4_14.INJECT1_0 = "NO";
    defparam phase_accum_add_4_14.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_12 (.A0(phase_inc_carrGen1[10]), .B0(phase_accum_adj_5658[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[11]), .B1(phase_accum_adj_5658[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15627), .COUT(n15628), .S0(n291), 
          .S1(n288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_12.INIT0 = 16'h666a;
    defparam phase_accum_add_4_12.INIT1 = 16'h666a;
    defparam phase_accum_add_4_12.INJECT1_0 = "NO";
    defparam phase_accum_add_4_12.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_10 (.A0(phase_inc_carrGen1[8]), .B0(phase_accum_adj_5658[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[9]), .B1(phase_accum_adj_5658[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15626), .COUT(n15627), .S0(n297), 
          .S1(n294));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_10.INIT0 = 16'h666a;
    defparam phase_accum_add_4_10.INIT1 = 16'h666a;
    defparam phase_accum_add_4_10.INJECT1_0 = "NO";
    defparam phase_accum_add_4_10.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_8 (.A0(phase_inc_carrGen1[6]), .B0(phase_accum_adj_5658[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[7]), .B1(phase_accum_adj_5658[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15625), .COUT(n15626), .S0(n303), 
          .S1(n300));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_8.INIT0 = 16'h666a;
    defparam phase_accum_add_4_8.INIT1 = 16'h666a;
    defparam phase_accum_add_4_8.INJECT1_0 = "NO";
    defparam phase_accum_add_4_8.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_6 (.A0(phase_inc_carrGen1[4]), .B0(phase_accum_adj_5658[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[5]), .B1(phase_accum_adj_5658[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15624), .COUT(n15625), .S0(n309), 
          .S1(n306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_6.INIT0 = 16'h666a;
    defparam phase_accum_add_4_6.INIT1 = 16'h666a;
    defparam phase_accum_add_4_6.INJECT1_0 = "NO";
    defparam phase_accum_add_4_6.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_4 (.A0(phase_inc_carrGen1[2]), .B0(phase_accum_adj_5658[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[3]), .B1(phase_accum_adj_5658[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15623), .COUT(n15624), .S0(n315), 
          .S1(n312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_4.INIT0 = 16'h666a;
    defparam phase_accum_add_4_4.INIT1 = 16'h666a;
    defparam phase_accum_add_4_4.INJECT1_0 = "NO";
    defparam phase_accum_add_4_4.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_2 (.A0(phase_inc_carrGen1[0]), .B0(phase_accum_adj_5658[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[1]), .B1(phase_accum_adj_5658[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15623), .S1(n318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_add_4_2.INIT0 = 16'h0008;
    defparam phase_accum_add_4_2.INIT1 = 16'h666a;
    defparam phase_accum_add_4_2.INJECT1_0 = "NO";
    defparam phase_accum_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_12 (.A0(counter[9]), .B0(DataInReg[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15621), .S1(cout_adj_4998));
    defparam _add_1_1649_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_12.INIT1 = 16'h0000;
    defparam _add_1_1649_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_10 (.A0(counter[7]), .B0(DataInReg[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(DataInReg[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15620), .COUT(n15621));
    defparam _add_1_1649_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_8 (.A0(counter[5]), .B0(DataInReg[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(DataInReg[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15619), .COUT(n15620));
    defparam _add_1_1649_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_6 (.A0(counter[3]), .B0(DataInReg[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(DataInReg[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15618), .COUT(n15619));
    defparam _add_1_1649_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_4 (.A0(counter[1]), .B0(DataInReg[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(DataInReg[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15617), .COUT(n15618));
    defparam _add_1_1649_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1649_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1649_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[0]), .B1(DataInReg[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15617));
    defparam _add_1_1649_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1649_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1649_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1649_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_13 (.A0(LOSine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15616), .S0(MixerOutSin_11__N_236[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1454_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_11 (.A0(LOSine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15615), .COUT(n15616), .S0(MixerOutSin_11__N_236[9]), 
          .S1(MixerOutSin_11__N_236[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_9 (.A0(LOSine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15614), .COUT(n15615), .S0(MixerOutSin_11__N_236[7]), 
          .S1(MixerOutSin_11__N_236[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_7 (.A0(LOSine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15613), .COUT(n15614), .S0(MixerOutSin_11__N_236[5]), 
          .S1(MixerOutSin_11__N_236[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_5 (.A0(LOSine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15612), .COUT(n15613), .S0(MixerOutSin_11__N_236[3]), 
          .S1(MixerOutSin_11__N_236[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_3 (.A0(LOSine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15611), .COUT(n15612), .S0(MixerOutSin_11__N_236[1]), 
          .S1(MixerOutSin_11__N_236[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1454_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1454_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_3.INJECT1_1 = "NO";
    LUT4 mux_325_i19_4_lut (.A(n11949), .B(n265), .C(n17625), .D(n2571), 
         .Z(n2352)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i19_4_lut.init = 16'hc0ca;
    CCU2C add_3639_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(ISquare[0]), 
          .A1(d_out_d_11__N_1892[17]), .B1(ISquare[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16366));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(58[15:27])
    defparam add_3639_1.INIT0 = 16'h000A;
    defparam add_3639_1.INIT1 = 16'h666a;
    defparam add_3639_1.INJECT1_0 = "NO";
    defparam add_3639_1.INJECT1_1 = "NO";
    LUT4 i3409_2_lut_2_lut (.A(o_Rx_Byte[3]), .B(n226_adj_5630), .Z(n2541)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3409_2_lut_2_lut.init = 16'hdddd;
    LUT4 i348_2_lut_rep_156_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(o_Rx_Byte[0]), 
         .C(n17634), .D(o_Rx_Byte[4]), .Z(n17625)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i348_2_lut_rep_156_4_lut_4_lut.init = 16'h4000;
    LUT4 i3341_3_lut_3_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(n193_adj_5619), 
         .C(n17633), .D(n12378), .Z(n2530)) /* synthesis lut_function=(A (B)+!A !(C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3341_3_lut_3_lut_4_lut_4_lut.init = 16'h8ddd;
    LUT4 i3338_3_lut_4_lut_3_lut (.A(o_Rx_Byte[3]), .B(n277_adj_5647), .C(n17630), 
         .Z(n2558)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3338_3_lut_4_lut_3_lut.init = 16'hd8d8;
    CCU2C add_3645_65 (.A0(phase_inc_carrGen[62]), .B0(n13169), .C0(n12146), 
          .D0(n3659), .A1(phase_inc_carrGen[63]), .B1(n13169), .C1(n12148), 
          .D1(n3659), .CIN(n16364), .S0(n137), .S1(n134));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_65.INIT0 = 16'h74b8;
    defparam add_3645_65.INIT1 = 16'h74b8;
    defparam add_3645_65.INJECT1_0 = "NO";
    defparam add_3645_65.INJECT1_1 = "NO";
    CCU2C add_3645_63 (.A0(phase_inc_carrGen[60]), .B0(n13169), .C0(n2310), 
          .D0(n3659), .A1(phase_inc_carrGen[61]), .B1(n13169), .C1(n12144), 
          .D1(n3659), .CIN(n16363), .COUT(n16364), .S0(n143), .S1(n140));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_63.INIT0 = 16'h74b8;
    defparam add_3645_63.INIT1 = 16'h74b8;
    defparam add_3645_63.INJECT1_0 = "NO";
    defparam add_3645_63.INJECT1_1 = "NO";
    LUT4 i2437_4_lut (.A(n262), .B(n256_adj_5640), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12138)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2437_4_lut.init = 16'hcac0;
    LUT4 mux_325_i17_4_lut (.A(n11945), .B(n271), .C(n17625), .D(n2571), 
         .Z(n2354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i17_4_lut.init = 16'hcfca;
    LUT4 i2246_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n286_adj_5650), 
         .Z(n11935)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2246_3_lut_4_lut.init = 16'hf707;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n17751), .B(o_Rx_Byte[2]), .C(n17633), 
         .D(n12378), .Z(n2636)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i3339_3_lut_3_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(n268_adj_5644), 
         .C(n17633), .D(n12378), .Z(n2555)) /* synthesis lut_function=(A (B)+!A !(C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3339_3_lut_3_lut_4_lut_4_lut.init = 16'h8ddd;
    LUT4 i2240_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n298_adj_5654), .Z(n11929)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2240_3_lut_4_lut.init = 16'hf808;
    CCU2C add_3645_61 (.A0(phase_inc_carrGen[58]), .B0(n13169), .C0(n2312), 
          .D0(n3659), .A1(phase_inc_carrGen[59]), .B1(n13169), .C1(n2311), 
          .D1(n3659), .CIN(n16362), .COUT(n16363), .S0(n149), .S1(n146));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_61.INIT0 = 16'h74b8;
    defparam add_3645_61.INIT1 = 16'h74b8;
    defparam add_3645_61.INJECT1_0 = "NO";
    defparam add_3645_61.INJECT1_1 = "NO";
    CCU2C add_3645_59 (.A0(phase_inc_carrGen[56]), .B0(n13169), .C0(n2314), 
          .D0(n3659), .A1(phase_inc_carrGen[57]), .B1(n13169), .C1(n2313), 
          .D1(n3659), .CIN(n16361), .COUT(n16362), .S0(n155), .S1(n152));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_59.INIT0 = 16'h74b8;
    defparam add_3645_59.INIT1 = 16'h74b8;
    defparam add_3645_59.INJECT1_0 = "NO";
    defparam add_3645_59.INJECT1_1 = "NO";
    LUT4 i3337_3_lut_3_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(n292_adj_5652), 
         .C(n17633), .D(n12378), .Z(n2563)) /* synthesis lut_function=(A (B)+!A !(C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3337_3_lut_3_lut_4_lut_4_lut.init = 16'h8ddd;
    LUT4 i3347_2_lut_2_lut (.A(o_Rx_Byte[3]), .B(n181_adj_5615), .Z(n2392)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3347_2_lut_2_lut.init = 16'hdddd;
    CCU2C add_3645_57 (.A0(phase_inc_carrGen[54]), .B0(n13169), .C0(n2316), 
          .D0(n3659), .A1(phase_inc_carrGen[55]), .B1(n13169), .C1(n2315), 
          .D1(n3659), .CIN(n16360), .COUT(n16361), .S0(n161), .S1(n158));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_57.INIT0 = 16'h74b8;
    defparam add_3645_57.INIT1 = 16'h74b8;
    defparam add_3645_57.INJECT1_0 = "NO";
    defparam add_3645_57.INJECT1_1 = "NO";
    LUT4 i3340_3_lut_3_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(n247_adj_5637), 
         .C(n17633), .D(n12378), .Z(n2548)) /* synthesis lut_function=(A (B)+!A !(C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3340_3_lut_3_lut_4_lut_4_lut.init = 16'h8ddd;
    CCU2C add_3645_55 (.A0(phase_inc_carrGen[52]), .B0(n13169), .C0(n12142), 
          .D0(n3659), .A1(phase_inc_carrGen[53]), .B1(n13169), .C1(n2317), 
          .D1(n3659), .CIN(n16359), .COUT(n16360), .S0(n167), .S1(n164));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_55.INIT0 = 16'h74b8;
    defparam add_3645_55.INIT1 = 16'h74b8;
    defparam add_3645_55.INJECT1_0 = "NO";
    defparam add_3645_55.INJECT1_1 = "NO";
    CCU2C add_3645_53 (.A0(phase_inc_carrGen[50]), .B0(n13169), .C0(n2320), 
          .D0(n3656), .A1(phase_inc_carrGen[51]), .B1(n13169), .C1(n2319), 
          .D1(n3659), .CIN(n16358), .COUT(n16359), .S0(n173), .S1(n170));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_53.INIT0 = 16'h74b8;
    defparam add_3645_53.INIT1 = 16'h74b8;
    defparam add_3645_53.INJECT1_0 = "NO";
    defparam add_3645_53.INJECT1_1 = "NO";
    LUT4 i2435_4_lut (.A(n268), .B(n262_adj_5642), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12136)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2435_4_lut.init = 16'hcac0;
    LUT4 i3262_4_lut (.A(n10_adj_4732), .B(n17098), .C(n16818), .D(n16812), 
         .Z(n12966)) /* synthesis lut_function=(A (B+(D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i3262_4_lut.init = 16'hfac8;
    CCU2C add_3645_51 (.A0(phase_inc_carrGen[48]), .B0(n13169), .C0(n2322), 
          .D0(n3656), .A1(phase_inc_carrGen[49]), .B1(n13169), .C1(n2321), 
          .D1(n3656), .CIN(n16357), .COUT(n16358), .S0(n179), .S1(n176));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_51.INIT0 = 16'h74b8;
    defparam add_3645_51.INIT1 = 16'h74b8;
    defparam add_3645_51.INJECT1_0 = "NO";
    defparam add_3645_51.INJECT1_1 = "NO";
    CCU2C add_3645_49 (.A0(phase_inc_carrGen[46]), .B0(n13169), .C0(n2324), 
          .D0(n11690), .A1(phase_inc_carrGen[47]), .B1(n13169), .C1(n2323), 
          .D1(n11690), .CIN(n16356), .COUT(n16357), .S0(n185), .S1(n182));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_49.INIT0 = 16'h74b8;
    defparam add_3645_49.INIT1 = 16'h74b8;
    defparam add_3645_49.INJECT1_0 = "NO";
    defparam add_3645_49.INJECT1_1 = "NO";
    CCU2C add_3645_47 (.A0(phase_inc_carrGen[44]), .B0(n13169), .C0(n2326), 
          .D0(n17622), .A1(phase_inc_carrGen[45]), .B1(n13169), .C1(n2325), 
          .D1(n3659), .CIN(n16355), .COUT(n16356), .S0(n191), .S1(n188));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_47.INIT0 = 16'h74b8;
    defparam add_3645_47.INIT1 = 16'h74b8;
    defparam add_3645_47.INJECT1_0 = "NO";
    defparam add_3645_47.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_30 (.A0(d1_adj_5667[63]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[64]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15284), .COUT(n15285), .S0(n102_adj_5445), 
          .S1(n99_adj_5444));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_28 (.A0(d1_adj_5667[61]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[62]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15283), .COUT(n15284), .S0(n108_adj_5447), 
          .S1(n105_adj_5446));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_26 (.A0(d1_adj_5667[59]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[60]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15282), .COUT(n15283), .S0(n114_adj_5449), 
          .S1(n111_adj_5448));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_24 (.A0(d1_adj_5667[57]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[58]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15281), .COUT(n15282), .S0(n120_adj_5451), 
          .S1(n117_adj_5450));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_22 (.A0(d1_adj_5667[55]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[56]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15280), .COUT(n15281), .S0(n126_adj_5453), 
          .S1(n123_adj_5452));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_20 (.A0(d1_adj_5667[53]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[54]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15279), .COUT(n15280), .S0(n132_adj_5455), 
          .S1(n129_adj_5454));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_18 (.A0(d1_adj_5667[51]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[52]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15278), .COUT(n15279), .S0(n138_adj_5457), 
          .S1(n135_adj_5456));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_16 (.A0(d1_adj_5667[49]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[50]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15277), .COUT(n15278), .S0(n144_adj_5459), 
          .S1(n141_adj_5458));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_14 (.A0(d1_adj_5667[47]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[48]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15276), .COUT(n15277), .S0(n150_adj_5461), 
          .S1(n147_adj_5460));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_12 (.A0(d1_adj_5667[45]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[46]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15275), .COUT(n15276), .S0(n156_adj_5463), 
          .S1(n153_adj_5462));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_10 (.A0(d1_adj_5667[43]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[44]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15274), .COUT(n15275), .S0(n162_adj_5465), 
          .S1(n159_adj_5464));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_8 (.A0(d1_adj_5667[41]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[42]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15273), .COUT(n15274), .S0(n168_adj_5467), 
          .S1(n165_adj_5466));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_6 (.A0(d1_adj_5667[39]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[40]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15272), .COUT(n15273), .S0(n174_adj_5469), 
          .S1(n171_adj_5468));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_4 (.A0(d1_adj_5667[37]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[38]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15271), .COUT(n15272), .S0(n180_adj_5471), 
          .S1(n177_adj_5470));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1565_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1_adj_5667[36]), .B1(MixerOutCos[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15271), .S1(n183_adj_5472));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1565_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1565_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1565_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_38 (.A0(d2[71]), .B0(d1[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15270), .S0(n78_adj_5180));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1553_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_36 (.A0(d2[69]), .B0(d1[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[70]), .B1(d1[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15269), .COUT(n15270), .S0(n84_adj_5182), .S1(n81_adj_5181));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_34 (.A0(d2[67]), .B0(d1[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[68]), .B1(d1[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15268), .COUT(n15269), .S0(n90_adj_5184), .S1(n87_adj_5183));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_32 (.A0(d2[65]), .B0(d1[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[66]), .B1(d1[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15267), .COUT(n15268), .S0(n96_adj_5186), .S1(n93_adj_5185));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_30 (.A0(d2[63]), .B0(d1[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[64]), .B1(d1[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15266), .COUT(n15267), .S0(n102_adj_5188), .S1(n99_adj_5187));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_28 (.A0(d2[61]), .B0(d1[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[62]), .B1(d1[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15265), .COUT(n15266), .S0(n108_adj_5190), .S1(n105_adj_5189));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_26 (.A0(d2[59]), .B0(d1[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[60]), .B1(d1[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15264), .COUT(n15265), .S0(n114_adj_5192), .S1(n111_adj_5191));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_24 (.A0(d2[57]), .B0(d1[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[58]), .B1(d1[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15263), .COUT(n15264), .S0(n120_adj_5194), .S1(n117_adj_5193));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_22 (.A0(d2[55]), .B0(d1[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[56]), .B1(d1[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15262), .COUT(n15263), .S0(n126_adj_5196), .S1(n123_adj_5195));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_20 (.A0(d2[53]), .B0(d1[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[54]), .B1(d1[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15261), .COUT(n15262), .S0(n132_adj_5198), .S1(n129_adj_5197));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_18 (.A0(d2[51]), .B0(d1[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[52]), .B1(d1[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15260), .COUT(n15261), .S0(n138_adj_5200), .S1(n135_adj_5199));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_16 (.A0(d2[49]), .B0(d1[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[50]), .B1(d1[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15259), .COUT(n15260), .S0(n144_adj_5202), .S1(n141_adj_5201));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_14 (.A0(d2[47]), .B0(d1[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[48]), .B1(d1[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15258), .COUT(n15259), .S0(n150_adj_5204), .S1(n147_adj_5203));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_12 (.A0(d2[45]), .B0(d1[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[46]), .B1(d1[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15257), .COUT(n15258), .S0(n156_adj_5206), .S1(n153_adj_5205));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_10 (.A0(d2[43]), .B0(d1[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[44]), .B1(d1[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15256), .COUT(n15257), .S0(n162_adj_5208), .S1(n159_adj_5207));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_8 (.A0(d2[41]), .B0(d1[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[42]), .B1(d1[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15255), .COUT(n15256), .S0(n168_adj_5210), .S1(n165_adj_5209));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_6 (.A0(d2[39]), .B0(d1[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[40]), .B1(d1[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15254), .COUT(n15255), .S0(n174_adj_5212), .S1(n171_adj_5211));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_4 (.A0(d2[37]), .B0(d1[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[38]), .B1(d1[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15253), .COUT(n15254), .S0(n180_adj_5214), .S1(n177_adj_5213));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[36]), .B1(d1[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15253), .S1(n183_adj_5215));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1553_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1553_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_38 (.A0(d_d8_adj_5677[35]), .B0(d8_adj_5676[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15252), .S0(d9_71__N_1675_adj_5702[35]), 
          .S1(cout_adj_5216));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1601_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_36 (.A0(d_d8_adj_5677[33]), .B0(d8_adj_5676[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[34]), .B1(d8_adj_5676[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15251), .COUT(n15252), .S0(d9_71__N_1675_adj_5702[33]), 
          .S1(d9_71__N_1675_adj_5702[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_34 (.A0(d_d8_adj_5677[31]), .B0(d8_adj_5676[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[32]), .B1(d8_adj_5676[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15250), .COUT(n15251), .S0(d9_71__N_1675_adj_5702[31]), 
          .S1(d9_71__N_1675_adj_5702[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_32 (.A0(d_d8_adj_5677[29]), .B0(d8_adj_5676[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[30]), .B1(d8_adj_5676[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15249), .COUT(n15250), .S0(d9_71__N_1675_adj_5702[29]), 
          .S1(d9_71__N_1675_adj_5702[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_30 (.A0(d_d8_adj_5677[27]), .B0(d8_adj_5676[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[28]), .B1(d8_adj_5676[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15248), .COUT(n15249), .S0(d9_71__N_1675_adj_5702[27]), 
          .S1(d9_71__N_1675_adj_5702[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_28 (.A0(d_d8_adj_5677[25]), .B0(d8_adj_5676[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[26]), .B1(d8_adj_5676[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15247), .COUT(n15248), .S0(d9_71__N_1675_adj_5702[25]), 
          .S1(d9_71__N_1675_adj_5702[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_26 (.A0(d_d8_adj_5677[23]), .B0(d8_adj_5676[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[24]), .B1(d8_adj_5676[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15246), .COUT(n15247), .S0(d9_71__N_1675_adj_5702[23]), 
          .S1(d9_71__N_1675_adj_5702[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_24 (.A0(d_d8_adj_5677[21]), .B0(d8_adj_5676[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[22]), .B1(d8_adj_5676[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15245), .COUT(n15246), .S0(d9_71__N_1675_adj_5702[21]), 
          .S1(d9_71__N_1675_adj_5702[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_22 (.A0(d_d8_adj_5677[19]), .B0(d8_adj_5676[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[20]), .B1(d8_adj_5676[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15244), .COUT(n15245), .S0(d9_71__N_1675_adj_5702[19]), 
          .S1(d9_71__N_1675_adj_5702[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_20 (.A0(d_d8_adj_5677[17]), .B0(d8_adj_5676[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[18]), .B1(d8_adj_5676[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15243), .COUT(n15244), .S0(d9_71__N_1675_adj_5702[17]), 
          .S1(d9_71__N_1675_adj_5702[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_18 (.A0(d_d8_adj_5677[15]), .B0(d8_adj_5676[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[16]), .B1(d8_adj_5676[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15242), .COUT(n15243), .S0(d9_71__N_1675_adj_5702[15]), 
          .S1(d9_71__N_1675_adj_5702[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_16 (.A0(d_d8_adj_5677[13]), .B0(d8_adj_5676[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[14]), .B1(d8_adj_5676[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15241), .COUT(n15242), .S0(d9_71__N_1675_adj_5702[13]), 
          .S1(d9_71__N_1675_adj_5702[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_14 (.A0(d_d8_adj_5677[11]), .B0(d8_adj_5676[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[12]), .B1(d8_adj_5676[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15240), .COUT(n15241), .S0(d9_71__N_1675_adj_5702[11]), 
          .S1(d9_71__N_1675_adj_5702[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_12 (.A0(d_d8_adj_5677[9]), .B0(d8_adj_5676[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[10]), .B1(d8_adj_5676[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15239), .COUT(n15240), .S0(d9_71__N_1675_adj_5702[9]), 
          .S1(d9_71__N_1675_adj_5702[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_10 (.A0(d_d8_adj_5677[7]), .B0(d8_adj_5676[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[8]), .B1(d8_adj_5676[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15238), .COUT(n15239), .S0(d9_71__N_1675_adj_5702[7]), 
          .S1(d9_71__N_1675_adj_5702[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_8 (.A0(d_d8_adj_5677[5]), .B0(d8_adj_5676[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[6]), .B1(d8_adj_5676[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15237), .COUT(n15238), .S0(d9_71__N_1675_adj_5702[5]), 
          .S1(d9_71__N_1675_adj_5702[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_6 (.A0(d_d8_adj_5677[3]), .B0(d8_adj_5676[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[4]), .B1(d8_adj_5676[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15236), .COUT(n15237), .S0(d9_71__N_1675_adj_5702[3]), 
          .S1(d9_71__N_1675_adj_5702[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_4 (.A0(d_d8_adj_5677[1]), .B0(d8_adj_5676[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5677[2]), .B1(d8_adj_5676[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15235), .COUT(n15236), .S0(d9_71__N_1675_adj_5702[1]), 
          .S1(d9_71__N_1675_adj_5702[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5677[0]), .B1(d8_adj_5676[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15235), .S1(d9_71__N_1675_adj_5702[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1601_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1601_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_38 (.A0(d1[71]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15234), .S0(n78_adj_5090));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1550_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_36 (.A0(d1[69]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[70]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15233), .COUT(n15234), .S0(n84_adj_5092), 
          .S1(n81_adj_5091));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_34 (.A0(d1[67]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[68]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15232), .COUT(n15233), .S0(n90_adj_5094), 
          .S1(n87_adj_5093));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_32 (.A0(d1[65]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[66]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15231), .COUT(n15232), .S0(n96_adj_5096), 
          .S1(n93_adj_5095));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_30 (.A0(d1[63]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[64]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15230), .COUT(n15231), .S0(n102_adj_5098), 
          .S1(n99_adj_5097));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_28 (.A0(d1[61]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[62]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15229), .COUT(n15230), .S0(n108_adj_5100), 
          .S1(n105_adj_5099));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_26 (.A0(d1[59]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[60]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15228), .COUT(n15229), .S0(n114_adj_5102), 
          .S1(n111_adj_5101));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_24 (.A0(d1[57]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[58]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15227), .COUT(n15228), .S0(n120_adj_5104), 
          .S1(n117_adj_5103));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_22 (.A0(d1[55]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[56]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15226), .COUT(n15227), .S0(n126_adj_5106), 
          .S1(n123_adj_5105));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_20 (.A0(d1[53]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[54]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15225), .COUT(n15226), .S0(n132_adj_5108), 
          .S1(n129_adj_5107));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_18 (.A0(d1[51]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[52]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15224), .COUT(n15225), .S0(n138_adj_5110), 
          .S1(n135_adj_5109));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_16 (.A0(d1[49]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[50]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15223), .COUT(n15224), .S0(n144_adj_5112), 
          .S1(n141_adj_5111));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_14 (.A0(d1[47]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[48]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15222), .COUT(n15223), .S0(n150_adj_5114), 
          .S1(n147_adj_5113));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_12 (.A0(d1[45]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[46]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15221), .COUT(n15222), .S0(n156_adj_5116), 
          .S1(n153_adj_5115));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_10 (.A0(d1[43]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[44]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15220), .COUT(n15221), .S0(n162_adj_5118), 
          .S1(n159_adj_5117));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_8 (.A0(d1[41]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[42]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15219), .COUT(n15220), .S0(n168_adj_5120), 
          .S1(n165_adj_5119));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_6 (.A0(d1[39]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[40]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15218), .COUT(n15219), .S0(n174_adj_5122), 
          .S1(n171_adj_5121));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_4 (.A0(d1[37]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[38]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15217), .COUT(n15218), .S0(n180_adj_5124), 
          .S1(n177_adj_5123));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[36]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15217), .S1(n183_adj_5125));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1550_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1550_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15216), .S0(cout_adj_5126));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1421_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1421_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_36 (.A0(d4[34]), .B0(d3[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[35]), .B1(d3[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15215), .COUT(n15216), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_34 (.A0(d4[32]), .B0(d3[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[33]), .B1(d3[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15214), .COUT(n15215), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_32 (.A0(d4[30]), .B0(d3[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[31]), .B1(d3[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15213), .COUT(n15214), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_30 (.A0(d4[28]), .B0(d3[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[29]), .B1(d3[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15212), .COUT(n15213), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_28 (.A0(d4[26]), .B0(d3[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[27]), .B1(d3[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15211), .COUT(n15212), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_26 (.A0(d4[24]), .B0(d3[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[25]), .B1(d3[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15210), .COUT(n15211), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_24 (.A0(d4[22]), .B0(d3[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[23]), .B1(d3[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15209), .COUT(n15210), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_22 (.A0(d4[20]), .B0(d3[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[21]), .B1(d3[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15208), .COUT(n15209), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_20 (.A0(d4[18]), .B0(d3[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[19]), .B1(d3[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15207), .COUT(n15208), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_18 (.A0(d4[16]), .B0(d3[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[17]), .B1(d3[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15206), .COUT(n15207), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_16 (.A0(d4[14]), .B0(d3[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[15]), .B1(d3[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15205), .COUT(n15206), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_14 (.A0(d4[12]), .B0(d3[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[13]), .B1(d3[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15204), .COUT(n15205), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_12 (.A0(d4[10]), .B0(d3[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[11]), .B1(d3[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15203), .COUT(n15204), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_10 (.A0(d4[8]), .B0(d3[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[9]), .B1(d3[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15202), .COUT(n15203), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_8 (.A0(d4[6]), .B0(d3[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[7]), .B1(d3[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15201), 
          .COUT(n15202), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_6 (.A0(d4[4]), .B0(d3[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[5]), .B1(d3[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15200), 
          .COUT(n15201), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_4 (.A0(d4[2]), .B0(d3[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[3]), .B1(d3[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15199), 
          .COUT(n15200), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_2 (.A0(d4[0]), .B0(d3[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[1]), .B1(d3[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15199), 
          .S1(d4_71__N_634[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1421_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1421_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_2.INJECT1_1 = "NO";
    LUT4 n17027_bdd_4_lut (.A(n17027), .B(n16930), .C(n17750), .D(n12378), 
         .Z(n2823)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n17027_bdd_4_lut.init = 16'hca00;
    CCU2C _add_1_1424_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15197), .S0(cout_adj_5127));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1424_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1424_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_36 (.A0(d5[34]), .B0(d4[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[35]), .B1(d4[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15196), .COUT(n15197), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_34 (.A0(d5[32]), .B0(d4[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[33]), .B1(d4[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15195), .COUT(n15196), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_32 (.A0(d5[30]), .B0(d4[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[31]), .B1(d4[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15194), .COUT(n15195), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_30 (.A0(d5[28]), .B0(d4[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[29]), .B1(d4[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15193), .COUT(n15194), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_28 (.A0(d5[26]), .B0(d4[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[27]), .B1(d4[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15192), .COUT(n15193), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_26 (.A0(d5[24]), .B0(d4[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[25]), .B1(d4[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15191), .COUT(n15192), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_24 (.A0(d5[22]), .B0(d4[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[23]), .B1(d4[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15190), .COUT(n15191), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_22 (.A0(d5[20]), .B0(d4[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[21]), .B1(d4[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15189), .COUT(n15190), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_20 (.A0(d5[18]), .B0(d4[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[19]), .B1(d4[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15188), .COUT(n15189), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_18 (.A0(d5[16]), .B0(d4[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[17]), .B1(d4[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15187), .COUT(n15188), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_16 (.A0(d5[14]), .B0(d4[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[15]), .B1(d4[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15186), .COUT(n15187), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_14 (.A0(d5[12]), .B0(d4[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[13]), .B1(d4[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15185), .COUT(n15186), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_12 (.A0(d5[10]), .B0(d4[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[11]), .B1(d4[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15184), .COUT(n15185), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_10 (.A0(d5[8]), .B0(d4[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[9]), .B1(d4[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15183), .COUT(n15184), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_8 (.A0(d5[6]), .B0(d4[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[7]), .B1(d4[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15182), 
          .COUT(n15183), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_6 (.A0(d5[4]), .B0(d4[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[5]), .B1(d4[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15181), 
          .COUT(n15182), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_4 (.A0(d5[2]), .B0(d4[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[3]), .B1(d4[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15180), 
          .COUT(n15181), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_2 (.A0(d5[0]), .B0(d4[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[1]), .B1(d4[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15180), 
          .S1(d5_71__N_706[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1424_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1424_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15178), .S0(cout_adj_5128));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1427_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1427_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_36 (.A0(d1_adj_5667[34]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[35]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15177), .COUT(n15178), .S0(d1_71__N_418_adj_5683[34]), 
          .S1(d1_71__N_418_adj_5683[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_34 (.A0(d1_adj_5667[32]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[33]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15176), .COUT(n15177), .S0(d1_71__N_418_adj_5683[32]), 
          .S1(d1_71__N_418_adj_5683[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_32 (.A0(d1_adj_5667[30]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[31]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15175), .COUT(n15176), .S0(d1_71__N_418_adj_5683[30]), 
          .S1(d1_71__N_418_adj_5683[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_30 (.A0(d1_adj_5667[28]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[29]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15174), .COUT(n15175), .S0(d1_71__N_418_adj_5683[28]), 
          .S1(d1_71__N_418_adj_5683[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_28 (.A0(d1_adj_5667[26]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[27]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15173), .COUT(n15174), .S0(d1_71__N_418_adj_5683[26]), 
          .S1(d1_71__N_418_adj_5683[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_26 (.A0(d1_adj_5667[24]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[25]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15172), .COUT(n15173), .S0(d1_71__N_418_adj_5683[24]), 
          .S1(d1_71__N_418_adj_5683[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_24 (.A0(d1_adj_5667[22]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[23]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15171), .COUT(n15172), .S0(d1_71__N_418_adj_5683[22]), 
          .S1(d1_71__N_418_adj_5683[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_22 (.A0(d1_adj_5667[20]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[21]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15170), .COUT(n15171), .S0(d1_71__N_418_adj_5683[20]), 
          .S1(d1_71__N_418_adj_5683[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_20 (.A0(d1_adj_5667[18]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[19]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15169), .COUT(n15170), .S0(d1_71__N_418_adj_5683[18]), 
          .S1(d1_71__N_418_adj_5683[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_18 (.A0(d1_adj_5667[16]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[17]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15168), .COUT(n15169), .S0(d1_71__N_418_adj_5683[16]), 
          .S1(d1_71__N_418_adj_5683[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_16 (.A0(d1_adj_5667[14]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[15]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15167), .COUT(n15168), .S0(d1_71__N_418_adj_5683[14]), 
          .S1(d1_71__N_418_adj_5683[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_14 (.A0(d1_adj_5667[12]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[13]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15166), .COUT(n15167), .S0(d1_71__N_418_adj_5683[12]), 
          .S1(d1_71__N_418_adj_5683[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_12 (.A0(d1_adj_5667[10]), .B0(MixerOutCos[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[11]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15165), .COUT(n15166), .S0(d1_71__N_418_adj_5683[10]), 
          .S1(d1_71__N_418_adj_5683[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_10 (.A0(d1_adj_5667[8]), .B0(MixerOutCos[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[9]), .B1(MixerOutCos[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15164), .COUT(n15165), .S0(d1_71__N_418_adj_5683[8]), 
          .S1(d1_71__N_418_adj_5683[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_8 (.A0(d1_adj_5667[6]), .B0(MixerOutCos[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[7]), .B1(MixerOutCos[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15163), .COUT(n15164), .S0(d1_71__N_418_adj_5683[6]), 
          .S1(d1_71__N_418_adj_5683[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_6 (.A0(d1_adj_5667[4]), .B0(MixerOutCos[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[5]), .B1(MixerOutCos[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15162), .COUT(n15163), .S0(d1_71__N_418_adj_5683[4]), 
          .S1(d1_71__N_418_adj_5683[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_4 (.A0(d1_adj_5667[2]), .B0(MixerOutCos[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[3]), .B1(MixerOutCos[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15161), .COUT(n15162), .S0(d1_71__N_418_adj_5683[2]), 
          .S1(d1_71__N_418_adj_5683[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1427_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_2 (.A0(d1_adj_5667[0]), .B0(MixerOutCos[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5667[1]), .B1(MixerOutCos[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15161), .S1(d1_71__N_418_adj_5683[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1427_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1427_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1427_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15159), .S0(cout));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1415_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1415_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_36 (.A0(d2[34]), .B0(d1[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[35]), .B1(d1[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15158), .COUT(n15159), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_34 (.A0(d2[32]), .B0(d1[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[33]), .B1(d1[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15157), .COUT(n15158), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_32 (.A0(d2[30]), .B0(d1[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[31]), .B1(d1[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15156), .COUT(n15157), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_30 (.A0(d2[28]), .B0(d1[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[29]), .B1(d1[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15155), .COUT(n15156), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_28 (.A0(d2[26]), .B0(d1[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[27]), .B1(d1[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15154), .COUT(n15155), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_26 (.A0(d2[24]), .B0(d1[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[25]), .B1(d1[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15153), .COUT(n15154), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_24 (.A0(d2[22]), .B0(d1[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[23]), .B1(d1[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15152), .COUT(n15153), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_22 (.A0(d2[20]), .B0(d1[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[21]), .B1(d1[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15151), .COUT(n15152), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_20 (.A0(d2[18]), .B0(d1[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[19]), .B1(d1[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15150), .COUT(n15151), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_18 (.A0(d2[16]), .B0(d1[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[17]), .B1(d1[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15149), .COUT(n15150), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_16 (.A0(d2[14]), .B0(d1[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[15]), .B1(d1[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15148), .COUT(n15149), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_14 (.A0(d2[12]), .B0(d1[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[13]), .B1(d1[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15147), .COUT(n15148), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_12 (.A0(d2[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[11]), .B1(d1[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15146), .COUT(n15147), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_10 (.A0(d2[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[9]), .B1(d1[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15145), .COUT(n15146), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_8 (.A0(d2[6]), .B0(d1[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[7]), .B1(d1[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15144), 
          .COUT(n15145), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_6 (.A0(d2[4]), .B0(d1[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[5]), .B1(d1[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15143), 
          .COUT(n15144), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_4 (.A0(d2[2]), .B0(d1[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[3]), .B1(d1[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15142), 
          .COUT(n15143), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_2 (.A0(d2[0]), .B0(d1[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[1]), .B1(d1[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15142), 
          .S1(d2_71__N_490[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1415_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1415_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15140), .S0(cout_adj_4999));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1652_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1652_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_36 (.A0(d1[34]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[35]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15139), .COUT(n15140), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_34 (.A0(d1[32]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[33]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15138), .COUT(n15139), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_32 (.A0(d1[30]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[31]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15137), .COUT(n15138), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_30 (.A0(d1[28]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[29]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15136), .COUT(n15137), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_28 (.A0(d1[26]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[27]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15135), .COUT(n15136), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_26 (.A0(d1[24]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[25]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15134), .COUT(n15135), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_24 (.A0(d1[22]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[23]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15133), .COUT(n15134), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_22 (.A0(d1[20]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[21]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15132), .COUT(n15133), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_20 (.A0(d1[18]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[19]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15131), .COUT(n15132), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_18 (.A0(d1[16]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[17]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15130), .COUT(n15131), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_16 (.A0(d1[14]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[15]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15129), .COUT(n15130), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_14 (.A0(d1[12]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[13]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15128), .COUT(n15129), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_12 (.A0(d1[10]), .B0(MixerOutSin[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[11]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15127), .COUT(n15128), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_10 (.A0(d1[8]), .B0(MixerOutSin[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[9]), .B1(MixerOutSin[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15126), .COUT(n15127), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_8 (.A0(d1[6]), .B0(MixerOutSin[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[7]), .B1(MixerOutSin[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15125), .COUT(n15126), .S0(d1_71__N_418[6]), 
          .S1(d1_71__N_418[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_6 (.A0(d1[4]), .B0(MixerOutSin[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[5]), .B1(MixerOutSin[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15124), .COUT(n15125), .S0(d1_71__N_418[4]), 
          .S1(d1_71__N_418[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_4 (.A0(d1[2]), .B0(MixerOutSin[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[3]), .B1(MixerOutSin[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15123), .COUT(n15124), .S0(d1_71__N_418[2]), 
          .S1(d1_71__N_418[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1652_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1652_add_4_2 (.A0(d1[0]), .B0(MixerOutSin[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[1]), .B1(MixerOutSin[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15123), .S1(d1_71__N_418[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1652_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1652_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1652_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1652_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15121), .S0(cout_adj_4837));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1418_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1418_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_36 (.A0(d3[34]), .B0(d2[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[35]), .B1(d2[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15120), .COUT(n15121), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_34 (.A0(d3[32]), .B0(d2[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[33]), .B1(d2[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15119), .COUT(n15120), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_32 (.A0(d3[30]), .B0(d2[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[31]), .B1(d2[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15118), .COUT(n15119), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_30 (.A0(d3[28]), .B0(d2[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[29]), .B1(d2[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15117), .COUT(n15118), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_28 (.A0(d3[26]), .B0(d2[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[27]), .B1(d2[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15116), .COUT(n15117), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_26 (.A0(d3[24]), .B0(d2[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[25]), .B1(d2[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15115), .COUT(n15116), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_24 (.A0(d3[22]), .B0(d2[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[23]), .B1(d2[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15114), .COUT(n15115), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_22 (.A0(d3[20]), .B0(d2[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[21]), .B1(d2[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15113), .COUT(n15114), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_20 (.A0(d3[18]), .B0(d2[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[19]), .B1(d2[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15112), .COUT(n15113), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_18 (.A0(d3[16]), .B0(d2[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[17]), .B1(d2[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15111), .COUT(n15112), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_16 (.A0(d3[14]), .B0(d2[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[15]), .B1(d2[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15110), .COUT(n15111), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_14 (.A0(d3[12]), .B0(d2[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[13]), .B1(d2[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15109), .COUT(n15110), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_12 (.A0(d3[10]), .B0(d2[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[11]), .B1(d2[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15108), .COUT(n15109), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_10 (.A0(d3[8]), .B0(d2[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[9]), .B1(d2[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15107), .COUT(n15108), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_8 (.A0(d3[6]), .B0(d2[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[7]), .B1(d2[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15106), 
          .COUT(n15107), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_6 (.A0(d3[4]), .B0(d2[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[5]), .B1(d2[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15105), 
          .COUT(n15106), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_4 (.A0(d3[2]), .B0(d2[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[3]), .B1(d2[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15104), 
          .COUT(n15105), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_2 (.A0(d3[0]), .B0(d2[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[1]), .B1(d2[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15104), 
          .S1(d3_71__N_562[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1418_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1418_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_38 (.A0(d3_adj_5669[71]), .B0(d2_adj_5668[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15102), .S0(n78_adj_4838));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1571_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_36 (.A0(d3_adj_5669[69]), .B0(d2_adj_5668[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[70]), .B1(d2_adj_5668[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15101), .COUT(n15102), .S0(n84_adj_4840), 
          .S1(n81_adj_4839));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_34 (.A0(d3_adj_5669[67]), .B0(d2_adj_5668[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[68]), .B1(d2_adj_5668[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15100), .COUT(n15101), .S0(n90_adj_4842), 
          .S1(n87_adj_4841));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_32 (.A0(d3_adj_5669[65]), .B0(d2_adj_5668[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[66]), .B1(d2_adj_5668[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15099), .COUT(n15100), .S0(n96_adj_4844), 
          .S1(n93_adj_4843));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_30 (.A0(d3_adj_5669[63]), .B0(d2_adj_5668[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[64]), .B1(d2_adj_5668[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15098), .COUT(n15099), .S0(n102_adj_4846), 
          .S1(n99_adj_4845));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_28 (.A0(d3_adj_5669[61]), .B0(d2_adj_5668[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[62]), .B1(d2_adj_5668[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15097), .COUT(n15098), .S0(n108_adj_4848), 
          .S1(n105_adj_4847));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_26 (.A0(d3_adj_5669[59]), .B0(d2_adj_5668[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[60]), .B1(d2_adj_5668[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15096), .COUT(n15097), .S0(n114_adj_4850), 
          .S1(n111_adj_4849));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_24 (.A0(d3_adj_5669[57]), .B0(d2_adj_5668[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[58]), .B1(d2_adj_5668[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15095), .COUT(n15096), .S0(n120_adj_4852), 
          .S1(n117_adj_4851));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_22 (.A0(d3_adj_5669[55]), .B0(d2_adj_5668[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[56]), .B1(d2_adj_5668[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15094), .COUT(n15095), .S0(n126_adj_4854), 
          .S1(n123_adj_4853));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_20 (.A0(d3_adj_5669[53]), .B0(d2_adj_5668[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[54]), .B1(d2_adj_5668[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15093), .COUT(n15094), .S0(n132_adj_4856), 
          .S1(n129_adj_4855));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_18 (.A0(d3_adj_5669[51]), .B0(d2_adj_5668[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[52]), .B1(d2_adj_5668[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15092), .COUT(n15093), .S0(n138_adj_4858), 
          .S1(n135_adj_4857));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_16 (.A0(d3_adj_5669[49]), .B0(d2_adj_5668[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[50]), .B1(d2_adj_5668[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15091), .COUT(n15092), .S0(n144_adj_4860), 
          .S1(n141_adj_4859));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_14 (.A0(d3_adj_5669[47]), .B0(d2_adj_5668[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[48]), .B1(d2_adj_5668[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15090), .COUT(n15091), .S0(n150_adj_4862), 
          .S1(n147_adj_4861));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_12 (.A0(d3_adj_5669[45]), .B0(d2_adj_5668[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[46]), .B1(d2_adj_5668[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15089), .COUT(n15090), .S0(n156_adj_4864), 
          .S1(n153_adj_4863));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_10 (.A0(d3_adj_5669[43]), .B0(d2_adj_5668[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[44]), .B1(d2_adj_5668[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15088), .COUT(n15089), .S0(n162_adj_4866), 
          .S1(n159_adj_4865));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_8 (.A0(d3_adj_5669[41]), .B0(d2_adj_5668[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[42]), .B1(d2_adj_5668[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15087), .COUT(n15088), .S0(n168_adj_4868), 
          .S1(n165_adj_4867));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_6 (.A0(d3_adj_5669[39]), .B0(d2_adj_5668[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[40]), .B1(d2_adj_5668[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15086), .COUT(n15087), .S0(n174_adj_4870), 
          .S1(n171_adj_4869));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1571_add_4_4 (.A0(d3_adj_5669[37]), .B0(d2_adj_5668[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[38]), .B1(d2_adj_5668[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15085), .COUT(n15086), .S0(n180_adj_4872), 
          .S1(n177_adj_4871));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1571_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_4.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i2 (.D(n315), .CK(clk_80mhz), .Q(phase_accum_adj_5658[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i3 (.D(n312), .CK(clk_80mhz), .Q(phase_accum_adj_5658[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i4 (.D(n309), .CK(clk_80mhz), .Q(phase_accum_adj_5658[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i5 (.D(n306), .CK(clk_80mhz), .Q(phase_accum_adj_5658[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i6 (.D(n303), .CK(clk_80mhz), .Q(phase_accum_adj_5658[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i7 (.D(n300), .CK(clk_80mhz), .Q(phase_accum_adj_5658[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i8 (.D(n297), .CK(clk_80mhz), .Q(phase_accum_adj_5658[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i9 (.D(n294), .CK(clk_80mhz), .Q(phase_accum_adj_5658[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i10 (.D(n291), .CK(clk_80mhz), .Q(phase_accum_adj_5658[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i11 (.D(n288), .CK(clk_80mhz), .Q(phase_accum_adj_5658[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i12 (.D(n285), .CK(clk_80mhz), .Q(phase_accum_adj_5658[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i13 (.D(n282), .CK(clk_80mhz), .Q(phase_accum_adj_5658[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i14 (.D(n279), .CK(clk_80mhz), .Q(phase_accum_adj_5658[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i15 (.D(n276), .CK(clk_80mhz), .Q(phase_accum_adj_5658[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i16 (.D(n273), .CK(clk_80mhz), .Q(phase_accum_adj_5658[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i17 (.D(n270), .CK(clk_80mhz), .Q(phase_accum_adj_5658[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i18 (.D(n267), .CK(clk_80mhz), .Q(phase_accum_adj_5658[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i19 (.D(n264), .CK(clk_80mhz), .Q(phase_accum_adj_5658[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i20 (.D(n261), .CK(clk_80mhz), .Q(phase_accum_adj_5658[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i21 (.D(n258), .CK(clk_80mhz), .Q(phase_accum_adj_5658[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i22 (.D(n255), .CK(clk_80mhz), .Q(phase_accum_adj_5658[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i23 (.D(n252), .CK(clk_80mhz), .Q(phase_accum_adj_5658[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i24 (.D(n249), .CK(clk_80mhz), .Q(phase_accum_adj_5658[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i25 (.D(n246), .CK(clk_80mhz), .Q(phase_accum_adj_5658[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i26 (.D(n243), .CK(clk_80mhz), .Q(phase_accum_adj_5658[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i27 (.D(n240), .CK(clk_80mhz), .Q(phase_accum_adj_5658[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i28 (.D(n237), .CK(clk_80mhz), .Q(phase_accum_adj_5658[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i29 (.D(n234), .CK(clk_80mhz), .Q(phase_accum_adj_5658[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i30 (.D(n231), .CK(clk_80mhz), .Q(phase_accum_adj_5658[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i31 (.D(n228), .CK(clk_80mhz), .Q(phase_accum_adj_5658[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i32 (.D(n225), .CK(clk_80mhz), .Q(phase_accum_adj_5658[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i33 (.D(n222), .CK(clk_80mhz), .Q(phase_accum_adj_5658[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i34 (.D(n219), .CK(clk_80mhz), .Q(phase_accum_adj_5658[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i35 (.D(n216), .CK(clk_80mhz), .Q(phase_accum_adj_5658[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i36 (.D(n213), .CK(clk_80mhz), .Q(phase_accum_adj_5658[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i37 (.D(n210), .CK(clk_80mhz), .Q(phase_accum_adj_5658[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i38 (.D(n207), .CK(clk_80mhz), .Q(phase_accum_adj_5658[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i39 (.D(n204), .CK(clk_80mhz), .Q(phase_accum_adj_5658[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i40 (.D(n201), .CK(clk_80mhz), .Q(phase_accum_adj_5658[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i41 (.D(n198), .CK(clk_80mhz), .Q(phase_accum_adj_5658[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i42 (.D(n195), .CK(clk_80mhz), .Q(phase_accum_adj_5658[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i43 (.D(n192), .CK(clk_80mhz), .Q(phase_accum_adj_5658[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i44 (.D(n189), .CK(clk_80mhz), .Q(phase_accum_adj_5658[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i45 (.D(n186), .CK(clk_80mhz), .Q(phase_accum_adj_5658[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i46 (.D(n183_adj_4521), .CK(clk_80mhz), .Q(phase_accum_adj_5658[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i47 (.D(n180_adj_4522), .CK(clk_80mhz), .Q(phase_accum_adj_5658[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i48 (.D(n177_adj_4523), .CK(clk_80mhz), .Q(phase_accum_adj_5658[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i49 (.D(n174_adj_4524), .CK(clk_80mhz), .Q(phase_accum_adj_5658[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i50 (.D(n171_adj_4525), .CK(clk_80mhz), .Q(phase_accum_adj_5658[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i51 (.D(n168_adj_4526), .CK(clk_80mhz), .Q(phase_accum_adj_5658[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i52 (.D(n165_adj_4527), .CK(clk_80mhz), .Q(phase_accum_adj_5658[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i53 (.D(n162_adj_4528), .CK(clk_80mhz), .Q(phase_accum_adj_5658[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i54 (.D(n159_adj_4529), .CK(clk_80mhz), .Q(phase_accum_adj_5658[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i55 (.D(n156_adj_4530), .CK(clk_80mhz), .Q(phase_accum_adj_5658[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i56 (.D(n153_adj_4531), .CK(clk_80mhz), .Q(phase_accum[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i57 (.D(n150_adj_4532), .CK(clk_80mhz), .Q(phase_accum[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i58 (.D(n147_adj_4533), .CK(clk_80mhz), .Q(phase_accum[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i59 (.D(n144_adj_4534), .CK(clk_80mhz), .Q(phase_accum[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i60 (.D(n141_adj_4535), .CK(clk_80mhz), .Q(phase_accum[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i61 (.D(n138_adj_4536), .CK(clk_80mhz), .Q(phase_accum[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i62 (.D(n135_adj_4537), .CK(clk_80mhz), .Q(phase_accum[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i63 (.D(n132_adj_4538), .CK(clk_80mhz), .Q(phase_accum[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(37[17:45])
    defparam phase_accum_e3_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_1571_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3_adj_5669[36]), .B1(d2_adj_5668[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15085), .S1(n183_adj_4873));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1571_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1571_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1571_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1571_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_61 (.A0(phase_inc_carrGen[63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15084), .S0(n124));
    defparam _add_1_1406_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_1406_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_59 (.A0(phase_inc_carrGen[61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15083), .COUT(n15084), .S0(n130_adj_5598), 
          .S1(n127));
    defparam _add_1_1406_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_57 (.A0(phase_inc_carrGen[59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15082), .COUT(n15083), .S0(n136_adj_5600), 
          .S1(n133_adj_5599));
    defparam _add_1_1406_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_55 (.A0(phase_inc_carrGen[57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15081), .COUT(n15082), .S0(n142_adj_5602), 
          .S1(n139_adj_5601));
    defparam _add_1_1406_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_53 (.A0(phase_inc_carrGen[55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15080), .COUT(n15081), .S0(n148_adj_5604), 
          .S1(n145_adj_5603));
    defparam _add_1_1406_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_51 (.A0(phase_inc_carrGen[53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15079), .COUT(n15080), .S0(n154_adj_5606), 
          .S1(n151_adj_5605));
    defparam _add_1_1406_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_49 (.A0(phase_inc_carrGen[51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15078), .COUT(n15079), .S0(n160_adj_5608), 
          .S1(n157_adj_5607));
    defparam _add_1_1406_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_47 (.A0(phase_inc_carrGen[49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15077), .COUT(n15078), .S0(n166_adj_5610), 
          .S1(n163_adj_5609));
    defparam _add_1_1406_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_45 (.A0(phase_inc_carrGen[47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15076), .COUT(n15077), .S0(n172_adj_5612), 
          .S1(n169_adj_5611));
    defparam _add_1_1406_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_43 (.A0(phase_inc_carrGen[45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15075), .COUT(n15076), .S0(n178_adj_5614), 
          .S1(n175_adj_5613));
    defparam _add_1_1406_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_41 (.A0(phase_inc_carrGen[43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15074), .COUT(n15075), .S0(n184_adj_5616), 
          .S1(n181_adj_5615));
    defparam _add_1_1406_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_39 (.A0(phase_inc_carrGen[41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15073), .COUT(n15074), .S0(n190_adj_5618), 
          .S1(n187_adj_5617));
    defparam _add_1_1406_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_37 (.A0(phase_inc_carrGen[39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15072), .COUT(n15073), .S0(n196_adj_5620), 
          .S1(n193_adj_5619));
    defparam _add_1_1406_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_35 (.A0(phase_inc_carrGen[37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15071), .COUT(n15072), .S0(n202_adj_5622), 
          .S1(n199_adj_5621));
    defparam _add_1_1406_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_33 (.A0(phase_inc_carrGen[35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15070), .COUT(n15071), .S0(n208_adj_5624), 
          .S1(n205_adj_5623));
    defparam _add_1_1406_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_31 (.A0(phase_inc_carrGen[33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15069), .COUT(n15070), .S0(n214_adj_5626), 
          .S1(n211_adj_5625));
    defparam _add_1_1406_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_29 (.A0(phase_inc_carrGen[31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15068), .COUT(n15069), .S0(n220_adj_5628), 
          .S1(n217_adj_5627));
    defparam _add_1_1406_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_27 (.A0(phase_inc_carrGen[29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15067), .COUT(n15068), .S0(n226_adj_5630), 
          .S1(n223_adj_5629));
    defparam _add_1_1406_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_25 (.A0(phase_inc_carrGen[27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15066), .COUT(n15067), .S0(n232_adj_5632), 
          .S1(n229_adj_5631));
    defparam _add_1_1406_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_23 (.A0(phase_inc_carrGen[25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15065), .COUT(n15066), .S0(n238_adj_5634), 
          .S1(n235_adj_5633));
    defparam _add_1_1406_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_21 (.A0(phase_inc_carrGen[23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15064), .COUT(n15065), .S0(n244_adj_5636), 
          .S1(n241_adj_5635));
    defparam _add_1_1406_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_19 (.A0(phase_inc_carrGen[21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15063), .COUT(n15064), .S0(n250_adj_5638), 
          .S1(n247_adj_5637));
    defparam _add_1_1406_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_17 (.A0(phase_inc_carrGen[19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15062), .COUT(n15063), .S0(n256_adj_5640), 
          .S1(n253_adj_5639));
    defparam _add_1_1406_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_15 (.A0(phase_inc_carrGen[17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15061), .COUT(n15062), .S0(n262_adj_5642), 
          .S1(n259_adj_5641));
    defparam _add_1_1406_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_13 (.A0(phase_inc_carrGen[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15060), .COUT(n15061), .S0(n268_adj_5644), 
          .S1(n265_adj_5643));
    defparam _add_1_1406_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_11 (.A0(phase_inc_carrGen[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15059), .COUT(n15060), .S0(n274_adj_5646), 
          .S1(n271_adj_5645));
    defparam _add_1_1406_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_9 (.A0(phase_inc_carrGen[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15058), .COUT(n15059), .S0(n280_adj_5648), 
          .S1(n277_adj_5647));
    defparam _add_1_1406_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_7 (.A0(phase_inc_carrGen[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15057), .COUT(n15058), .S0(n286_adj_5650), 
          .S1(n283_adj_5649));
    defparam _add_1_1406_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_5 (.A0(phase_inc_carrGen[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15056), .COUT(n15057), .S0(n292_adj_5652), 
          .S1(n289_adj_5651));
    defparam _add_1_1406_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_1406_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_3 (.A0(phase_inc_carrGen[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15055), .COUT(n15056), .S0(n298_adj_5654), 
          .S1(n295_adj_5653));
    defparam _add_1_1406_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1406_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1406_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15055), .S1(n301_adj_5655));
    defparam _add_1_1406_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1406_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1406_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_38 (.A0(d_d7_adj_5675[35]), .B0(d7_adj_5674[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15054), .S0(d8_71__N_1603_adj_5701[35]), 
          .S1(cout_adj_5254));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1604_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_36 (.A0(d_d7_adj_5675[33]), .B0(d7_adj_5674[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[34]), .B1(d7_adj_5674[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15053), .COUT(n15054), .S0(d8_71__N_1603_adj_5701[33]), 
          .S1(d8_71__N_1603_adj_5701[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_34 (.A0(d_d7_adj_5675[31]), .B0(d7_adj_5674[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[32]), .B1(d7_adj_5674[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15052), .COUT(n15053), .S0(d8_71__N_1603_adj_5701[31]), 
          .S1(d8_71__N_1603_adj_5701[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_32 (.A0(d_d7_adj_5675[29]), .B0(d7_adj_5674[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[30]), .B1(d7_adj_5674[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15051), .COUT(n15052), .S0(d8_71__N_1603_adj_5701[29]), 
          .S1(d8_71__N_1603_adj_5701[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_30 (.A0(d_d7_adj_5675[27]), .B0(d7_adj_5674[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[28]), .B1(d7_adj_5674[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15050), .COUT(n15051), .S0(d8_71__N_1603_adj_5701[27]), 
          .S1(d8_71__N_1603_adj_5701[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_28 (.A0(d_d7_adj_5675[25]), .B0(d7_adj_5674[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[26]), .B1(d7_adj_5674[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15049), .COUT(n15050), .S0(d8_71__N_1603_adj_5701[25]), 
          .S1(d8_71__N_1603_adj_5701[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_26 (.A0(d_d7_adj_5675[23]), .B0(d7_adj_5674[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[24]), .B1(d7_adj_5674[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15048), .COUT(n15049), .S0(d8_71__N_1603_adj_5701[23]), 
          .S1(d8_71__N_1603_adj_5701[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_24 (.A0(d_d7_adj_5675[21]), .B0(d7_adj_5674[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[22]), .B1(d7_adj_5674[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15047), .COUT(n15048), .S0(d8_71__N_1603_adj_5701[21]), 
          .S1(d8_71__N_1603_adj_5701[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_22 (.A0(d_d7_adj_5675[19]), .B0(d7_adj_5674[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[20]), .B1(d7_adj_5674[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15046), .COUT(n15047), .S0(d8_71__N_1603_adj_5701[19]), 
          .S1(d8_71__N_1603_adj_5701[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_20 (.A0(d_d7_adj_5675[17]), .B0(d7_adj_5674[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[18]), .B1(d7_adj_5674[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15045), .COUT(n15046), .S0(d8_71__N_1603_adj_5701[17]), 
          .S1(d8_71__N_1603_adj_5701[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_18 (.A0(d_d7_adj_5675[15]), .B0(d7_adj_5674[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[16]), .B1(d7_adj_5674[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15044), .COUT(n15045), .S0(d8_71__N_1603_adj_5701[15]), 
          .S1(d8_71__N_1603_adj_5701[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_16 (.A0(d_d7_adj_5675[13]), .B0(d7_adj_5674[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[14]), .B1(d7_adj_5674[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15043), .COUT(n15044), .S0(d8_71__N_1603_adj_5701[13]), 
          .S1(d8_71__N_1603_adj_5701[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_14 (.A0(d_d7_adj_5675[11]), .B0(d7_adj_5674[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[12]), .B1(d7_adj_5674[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15042), .COUT(n15043), .S0(d8_71__N_1603_adj_5701[11]), 
          .S1(d8_71__N_1603_adj_5701[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_12 (.A0(d_d7_adj_5675[9]), .B0(d7_adj_5674[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[10]), .B1(d7_adj_5674[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15041), .COUT(n15042), .S0(d8_71__N_1603_adj_5701[9]), 
          .S1(d8_71__N_1603_adj_5701[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_10 (.A0(d_d7_adj_5675[7]), .B0(d7_adj_5674[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[8]), .B1(d7_adj_5674[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15040), .COUT(n15041), .S0(d8_71__N_1603_adj_5701[7]), 
          .S1(d8_71__N_1603_adj_5701[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_8 (.A0(d_d7_adj_5675[5]), .B0(d7_adj_5674[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[6]), .B1(d7_adj_5674[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15039), .COUT(n15040), .S0(d8_71__N_1603_adj_5701[5]), 
          .S1(d8_71__N_1603_adj_5701[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_6 (.A0(d_d7_adj_5675[3]), .B0(d7_adj_5674[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[4]), .B1(d7_adj_5674[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15038), .COUT(n15039), .S0(d8_71__N_1603_adj_5701[3]), 
          .S1(d8_71__N_1603_adj_5701[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_4 (.A0(d_d7_adj_5675[1]), .B0(d7_adj_5674[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[2]), .B1(d7_adj_5674[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15037), .COUT(n15038), .S0(d8_71__N_1603_adj_5701[1]), 
          .S1(d8_71__N_1603_adj_5701[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1604_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5675[0]), .B1(d7_adj_5674[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15037), .S1(d8_71__N_1603_adj_5701[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1604_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1604_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1604_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_38 (.A0(d_d8[35]), .B0(d8[35]), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15036), 
          .S0(d9_71__N_1675[35]), .S1(cout_adj_5000));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_36 (.A0(d_d8[33]), .B0(d8[33]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[34]), .B1(d8[34]), .C1(GND_net), .D1(VCC_net), .CIN(n15035), 
          .COUT(n15036), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_34 (.A0(d_d8[31]), .B0(d8[31]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[32]), .B1(d8[32]), .C1(GND_net), .D1(VCC_net), .CIN(n15034), 
          .COUT(n15035), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_32 (.A0(d_d8[29]), .B0(d8[29]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[30]), .B1(d8[30]), .C1(GND_net), .D1(VCC_net), .CIN(n15033), 
          .COUT(n15034), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_30 (.A0(d_d8[27]), .B0(d8[27]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[28]), .B1(d8[28]), .C1(GND_net), .D1(VCC_net), .CIN(n15032), 
          .COUT(n15033), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(d_d8[25]), .B0(d8[25]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[26]), .B1(d8[26]), .C1(GND_net), .D1(VCC_net), .CIN(n15031), 
          .COUT(n15032), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(d_d8[23]), .B0(d8[23]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[24]), .B1(d8[24]), .C1(GND_net), .D1(VCC_net), .CIN(n15030), 
          .COUT(n15031), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_24 (.A0(d_d8[21]), .B0(d8[21]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[22]), .B1(d8[22]), .C1(GND_net), .D1(VCC_net), .CIN(n15029), 
          .COUT(n15030), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_22 (.A0(d_d8[19]), .B0(d8[19]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[20]), .B1(d8[20]), .C1(GND_net), .D1(VCC_net), .CIN(n15028), 
          .COUT(n15029), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_20 (.A0(d_d8[17]), .B0(d8[17]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[18]), .B1(d8[18]), .C1(GND_net), .D1(VCC_net), .CIN(n15027), 
          .COUT(n15028), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_18 (.A0(d_d8[15]), .B0(d8[15]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[16]), .B1(d8[16]), .C1(GND_net), .D1(VCC_net), .CIN(n15026), 
          .COUT(n15027), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_16 (.A0(d_d8[13]), .B0(d8[13]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[14]), .B1(d8[14]), .C1(GND_net), .D1(VCC_net), .CIN(n15025), 
          .COUT(n15026), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_14 (.A0(d_d8[11]), .B0(d8[11]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[12]), .B1(d8[12]), .C1(GND_net), .D1(VCC_net), .CIN(n15024), 
          .COUT(n15025), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_12 (.A0(d_d8[9]), .B0(d8[9]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[10]), .B1(d8[10]), .C1(GND_net), .D1(VCC_net), .CIN(n15023), 
          .COUT(n15024), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_10 (.A0(d_d8[7]), .B0(d8[7]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[8]), .B1(d8[8]), .C1(GND_net), .D1(VCC_net), .CIN(n15022), 
          .COUT(n15023), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_8 (.A0(d_d8[5]), .B0(d8[5]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[6]), .B1(d8[6]), .C1(GND_net), .D1(VCC_net), .CIN(n15021), 
          .COUT(n15022), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_6 (.A0(d_d8[3]), .B0(d8[3]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[4]), .B1(d8[4]), .C1(GND_net), .D1(VCC_net), .CIN(n15020), 
          .COUT(n15021), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_4 (.A0(d_d8[1]), .B0(d8[1]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[2]), .B1(d8[2]), .C1(GND_net), .D1(VCC_net), .CIN(n15019), 
          .COUT(n15020), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[0]), .B1(d8[0]), .C1(GND_net), .D1(VCC_net), .COUT(n15019), 
          .S1(d9_71__N_1675[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_37 (.A0(d_d9_adj_5679[71]), .B0(d9_adj_5678[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15018), .S0(n76_adj_5521));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1469_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_35 (.A0(d_d9_adj_5679[69]), .B0(d9_adj_5678[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[70]), .B1(d9_adj_5678[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15017), .COUT(n15018), .S0(n82_adj_5523), 
          .S1(n79_adj_5522));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_33 (.A0(d_d9_adj_5679[67]), .B0(d9_adj_5678[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[68]), .B1(d9_adj_5678[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15016), .COUT(n15017), .S0(n88_adj_5525), 
          .S1(n85_adj_5524));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_31 (.A0(d_d9_adj_5679[65]), .B0(d9_adj_5678[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[66]), .B1(d9_adj_5678[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15015), .COUT(n15016), .S0(n94_adj_5527), 
          .S1(n91_adj_5526));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_29 (.A0(d_d9_adj_5679[63]), .B0(d9_adj_5678[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[64]), .B1(d9_adj_5678[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15014), .COUT(n15015), .S0(n100_adj_5529), 
          .S1(n97_adj_5528));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_27 (.A0(d_d9_adj_5679[61]), .B0(d9_adj_5678[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[62]), .B1(d9_adj_5678[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15013), .COUT(n15014), .S0(n106_adj_5531), 
          .S1(n103_adj_5530));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_25 (.A0(d_d9_adj_5679[59]), .B0(d9_adj_5678[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[60]), .B1(d9_adj_5678[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15012), .COUT(n15013), .S0(n112_adj_5533), 
          .S1(n109_adj_5532));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_23 (.A0(d_d9_adj_5679[57]), .B0(d9_adj_5678[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[58]), .B1(d9_adj_5678[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15011), .COUT(n15012), .S0(n118_adj_5535), 
          .S1(n115_adj_5534));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_21 (.A0(d_d9_adj_5679[55]), .B0(d9_adj_5678[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[56]), .B1(d9_adj_5678[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15010), .COUT(n15011));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_19 (.A0(d_d9_adj_5679[53]), .B0(d9_adj_5678[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[54]), .B1(d9_adj_5678[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15009), .COUT(n15010));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_17 (.A0(d_d9_adj_5679[51]), .B0(d9_adj_5678[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[52]), .B1(d9_adj_5678[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15008), .COUT(n15009));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_15 (.A0(d_d9_adj_5679[49]), .B0(d9_adj_5678[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[50]), .B1(d9_adj_5678[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15007), .COUT(n15008));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_13 (.A0(d_d9_adj_5679[47]), .B0(d9_adj_5678[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[48]), .B1(d9_adj_5678[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15006), .COUT(n15007));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_11 (.A0(d_d9_adj_5679[45]), .B0(d9_adj_5678[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[46]), .B1(d9_adj_5678[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15005), .COUT(n15006));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_9 (.A0(d_d9_adj_5679[43]), .B0(d9_adj_5678[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[44]), .B1(d9_adj_5678[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15004), .COUT(n15005));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_7 (.A0(d_d9_adj_5679[41]), .B0(d9_adj_5678[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[42]), .B1(d9_adj_5678[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15003), .COUT(n15004));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_5 (.A0(d_d9_adj_5679[39]), .B0(d9_adj_5678[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[40]), .B1(d9_adj_5678[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15002), .COUT(n15003));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_3 (.A0(d_d9_adj_5679[37]), .B0(d9_adj_5678[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[38]), .B1(d9_adj_5678[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15001), .COUT(n15002));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5679[36]), .B1(d9_adj_5678[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15001));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1469_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1469_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_38 (.A0(d_d9_adj_5679[71]), .B0(d9_adj_5678[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15000), .S0(n78_adj_4874));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1634_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_36 (.A0(d_d9_adj_5679[69]), .B0(d9_adj_5678[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[70]), .B1(d9_adj_5678[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14999), .COUT(n15000), .S0(n84_adj_4876), 
          .S1(n81_adj_4875));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_34 (.A0(d_d9_adj_5679[67]), .B0(d9_adj_5678[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[68]), .B1(d9_adj_5678[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14998), .COUT(n14999), .S0(n90_adj_4878), 
          .S1(n87_adj_4877));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_32 (.A0(d_d9_adj_5679[65]), .B0(d9_adj_5678[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[66]), .B1(d9_adj_5678[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14997), .COUT(n14998), .S0(n96_adj_4880), 
          .S1(n93_adj_4879));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_30 (.A0(d_d9_adj_5679[63]), .B0(d9_adj_5678[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[64]), .B1(d9_adj_5678[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14996), .COUT(n14997), .S0(n102_adj_4882), 
          .S1(n99_adj_4881));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_28 (.A0(d_d9_adj_5679[61]), .B0(d9_adj_5678[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[62]), .B1(d9_adj_5678[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14995), .COUT(n14996), .S0(n108_adj_4884), 
          .S1(n105_adj_4883));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_26 (.A0(d_d9_adj_5679[59]), .B0(d9_adj_5678[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[60]), .B1(d9_adj_5678[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14994), .COUT(n14995), .S0(n114_adj_4886), 
          .S1(n111_adj_4885));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_24 (.A0(d_d9_adj_5679[57]), .B0(d9_adj_5678[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[58]), .B1(d9_adj_5678[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14993), .COUT(n14994), .S0(n120_adj_4888), 
          .S1(n117_adj_4887));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_22 (.A0(d_d9_adj_5679[55]), .B0(d9_adj_5678[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[56]), .B1(d9_adj_5678[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14992), .COUT(n14993));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_20 (.A0(d_d9_adj_5679[53]), .B0(d9_adj_5678[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[54]), .B1(d9_adj_5678[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14991), .COUT(n14992));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_18 (.A0(d_d9_adj_5679[51]), .B0(d9_adj_5678[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[52]), .B1(d9_adj_5678[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14990), .COUT(n14991));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_16 (.A0(d_d9_adj_5679[49]), .B0(d9_adj_5678[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[50]), .B1(d9_adj_5678[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14989), .COUT(n14990));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_14 (.A0(d_d9_adj_5679[47]), .B0(d9_adj_5678[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[48]), .B1(d9_adj_5678[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14988), .COUT(n14989));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_12 (.A0(d_d9_adj_5679[45]), .B0(d9_adj_5678[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[46]), .B1(d9_adj_5678[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14987), .COUT(n14988));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_10 (.A0(d_d9_adj_5679[43]), .B0(d9_adj_5678[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[44]), .B1(d9_adj_5678[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14986), .COUT(n14987));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_8 (.A0(d_d9_adj_5679[41]), .B0(d9_adj_5678[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[42]), .B1(d9_adj_5678[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14985), .COUT(n14986));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_6 (.A0(d_d9_adj_5679[39]), .B0(d9_adj_5678[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[40]), .B1(d9_adj_5678[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14984), .COUT(n14985));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_4 (.A0(d_d9_adj_5679[37]), .B0(d9_adj_5678[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5679[38]), .B1(d9_adj_5678[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14983), .COUT(n14984));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1634_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1634_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5679[36]), .B1(d9_adj_5678[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14983));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1634_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1634_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1634_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1634_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_38 (.A0(d_d8[71]), .B0(d8[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14982), .S0(n78_adj_5001));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1580_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_36 (.A0(d_d8[69]), .B0(d8[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[70]), .B1(d8[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14981), .COUT(n14982), .S0(n84_adj_5003), .S1(n81_adj_5002));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_34 (.A0(d_d8[67]), .B0(d8[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[68]), .B1(d8[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14980), .COUT(n14981), .S0(n90_adj_5005), .S1(n87_adj_5004));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_32 (.A0(d_d8[65]), .B0(d8[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[66]), .B1(d8[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14979), .COUT(n14980), .S0(n96_adj_5007), .S1(n93_adj_5006));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_30 (.A0(d_d8[63]), .B0(d8[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[64]), .B1(d8[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14978), .COUT(n14979), .S0(n102_adj_5009), .S1(n99_adj_5008));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_28 (.A0(d_d8[61]), .B0(d8[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[62]), .B1(d8[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14977), .COUT(n14978), .S0(n108_adj_5011), .S1(n105_adj_5010));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_26 (.A0(d_d8[59]), .B0(d8[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[60]), .B1(d8[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14976), .COUT(n14977), .S0(n114_adj_5013), .S1(n111_adj_5012));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_24 (.A0(d_d8[57]), .B0(d8[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[58]), .B1(d8[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14975), .COUT(n14976), .S0(n120_adj_5015), .S1(n117_adj_5014));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_22 (.A0(d_d8[55]), .B0(d8[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[56]), .B1(d8[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14974), .COUT(n14975), .S0(n126_adj_5017), .S1(n123_adj_5016));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_20 (.A0(d_d8[53]), .B0(d8[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[54]), .B1(d8[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14973), .COUT(n14974), .S0(n132_adj_5019), .S1(n129_adj_5018));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_18 (.A0(d_d8[51]), .B0(d8[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[52]), .B1(d8[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14972), .COUT(n14973), .S0(n138_adj_5021), .S1(n135_adj_5020));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_16 (.A0(d_d8[49]), .B0(d8[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[50]), .B1(d8[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14971), .COUT(n14972), .S0(n144_adj_5023), .S1(n141_adj_5022));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_14 (.A0(d_d8[47]), .B0(d8[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[48]), .B1(d8[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14970), .COUT(n14971), .S0(n150_adj_5025), .S1(n147_adj_5024));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_12 (.A0(d_d8[45]), .B0(d8[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[46]), .B1(d8[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14969), .COUT(n14970), .S0(n156_adj_5027), .S1(n153_adj_5026));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_10 (.A0(d_d8[43]), .B0(d8[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[44]), .B1(d8[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14968), .COUT(n14969), .S0(n162_adj_5029), .S1(n159_adj_5028));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_8 (.A0(d_d8[41]), .B0(d8[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[42]), .B1(d8[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14967), .COUT(n14968), .S0(n168_adj_5031), .S1(n165_adj_5030));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_6 (.A0(d_d8[39]), .B0(d8[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[40]), .B1(d8[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14966), .COUT(n14967), .S0(n174_adj_5033), .S1(n171_adj_5032));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_4 (.A0(d_d8[37]), .B0(d8[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[38]), .B1(d8[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14965), .COUT(n14966), .S0(n180_adj_5035), .S1(n177_adj_5034));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[36]), .B1(d8[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n14965), .S1(n183_adj_5036));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam _add_1_1580_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1580_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14964), .S0(n36_adj_5129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1430_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14963), .COUT(n14964), .S0(n42), .S1(n39));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14962), .COUT(n14963), .S0(n48), .S1(n45));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14961), .COUT(n14962), .S0(n54), .S1(n51));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14960), .COUT(n14961), .S0(n60), .S1(n57));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14959), .COUT(n14960), .S0(n66_adj_5131), .S1(n63_adj_5130));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14958), .COUT(n14959), .S0(n72), .S1(n69));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14957), .COUT(n14958), .S0(n78_adj_5132), .S1(n75));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1430_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1430_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n14957), .S1(n81_adj_5133));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(87[24:37])
    defparam _add_1_1430_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1430_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1430_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_37 (.A0(d1[70]), .B0(cout), .C0(n81_adj_5181), 
          .D0(d2[70]), .A1(d1[71]), .B1(cout), .C1(n78_adj_5180), .D1(d2[71]), 
          .CIN(n14955), .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_35 (.A0(d1[68]), .B0(cout), .C0(n87_adj_5183), 
          .D0(d2[68]), .A1(d1[69]), .B1(cout), .C1(n84_adj_5182), .D1(d2[69]), 
          .CIN(n14954), .COUT(n14955), .S0(d2_71__N_490[68]), .S1(d2_71__N_490[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_33 (.A0(d1[66]), .B0(cout), .C0(n93_adj_5185), 
          .D0(d2[66]), .A1(d1[67]), .B1(cout), .C1(n90_adj_5184), .D1(d2[67]), 
          .CIN(n14953), .COUT(n14954), .S0(d2_71__N_490[66]), .S1(d2_71__N_490[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_31 (.A0(d1[64]), .B0(cout), .C0(n99_adj_5187), 
          .D0(d2[64]), .A1(d1[65]), .B1(cout), .C1(n96_adj_5186), .D1(d2[65]), 
          .CIN(n14952), .COUT(n14953), .S0(d2_71__N_490[64]), .S1(d2_71__N_490[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_29 (.A0(d1[62]), .B0(cout), .C0(n105_adj_5189), 
          .D0(d2[62]), .A1(d1[63]), .B1(cout), .C1(n102_adj_5188), .D1(d2[63]), 
          .CIN(n14951), .COUT(n14952), .S0(d2_71__N_490[62]), .S1(d2_71__N_490[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_27 (.A0(d1[60]), .B0(cout), .C0(n111_adj_5191), 
          .D0(d2[60]), .A1(d1[61]), .B1(cout), .C1(n108_adj_5190), .D1(d2[61]), 
          .CIN(n14950), .COUT(n14951), .S0(d2_71__N_490[60]), .S1(d2_71__N_490[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_25 (.A0(d1[58]), .B0(cout), .C0(n117_adj_5193), 
          .D0(d2[58]), .A1(d1[59]), .B1(cout), .C1(n114_adj_5192), .D1(d2[59]), 
          .CIN(n14949), .COUT(n14950), .S0(d2_71__N_490[58]), .S1(d2_71__N_490[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_23 (.A0(d1[56]), .B0(cout), .C0(n123_adj_5195), 
          .D0(d2[56]), .A1(d1[57]), .B1(cout), .C1(n120_adj_5194), .D1(d2[57]), 
          .CIN(n14948), .COUT(n14949), .S0(d2_71__N_490[56]), .S1(d2_71__N_490[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_21 (.A0(d1[54]), .B0(cout), .C0(n129_adj_5197), 
          .D0(d2[54]), .A1(d1[55]), .B1(cout), .C1(n126_adj_5196), .D1(d2[55]), 
          .CIN(n14947), .COUT(n14948), .S0(d2_71__N_490[54]), .S1(d2_71__N_490[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_19 (.A0(d1[52]), .B0(cout), .C0(n135_adj_5199), 
          .D0(d2[52]), .A1(d1[53]), .B1(cout), .C1(n132_adj_5198), .D1(d2[53]), 
          .CIN(n14946), .COUT(n14947), .S0(d2_71__N_490[52]), .S1(d2_71__N_490[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_17 (.A0(d1[50]), .B0(cout), .C0(n141_adj_5201), 
          .D0(d2[50]), .A1(d1[51]), .B1(cout), .C1(n138_adj_5200), .D1(d2[51]), 
          .CIN(n14945), .COUT(n14946), .S0(d2_71__N_490[50]), .S1(d2_71__N_490[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_15 (.A0(d1[48]), .B0(cout), .C0(n147_adj_5203), 
          .D0(d2[48]), .A1(d1[49]), .B1(cout), .C1(n144_adj_5202), .D1(d2[49]), 
          .CIN(n14944), .COUT(n14945), .S0(d2_71__N_490[48]), .S1(d2_71__N_490[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_13 (.A0(d1[46]), .B0(cout), .C0(n153_adj_5205), 
          .D0(d2[46]), .A1(d1[47]), .B1(cout), .C1(n150_adj_5204), .D1(d2[47]), 
          .CIN(n14943), .COUT(n14944), .S0(d2_71__N_490[46]), .S1(d2_71__N_490[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_11 (.A0(d1[44]), .B0(cout), .C0(n159_adj_5207), 
          .D0(d2[44]), .A1(d1[45]), .B1(cout), .C1(n156_adj_5206), .D1(d2[45]), 
          .CIN(n14942), .COUT(n14943), .S0(d2_71__N_490[44]), .S1(d2_71__N_490[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_9 (.A0(d1[42]), .B0(cout), .C0(n165_adj_5209), 
          .D0(d2[42]), .A1(d1[43]), .B1(cout), .C1(n162_adj_5208), .D1(d2[43]), 
          .CIN(n14941), .COUT(n14942), .S0(d2_71__N_490[42]), .S1(d2_71__N_490[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_7 (.A0(d1[40]), .B0(cout), .C0(n171_adj_5211), 
          .D0(d2[40]), .A1(d1[41]), .B1(cout), .C1(n168_adj_5210), .D1(d2[41]), 
          .CIN(n14940), .COUT(n14941), .S0(d2_71__N_490[40]), .S1(d2_71__N_490[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_5 (.A0(d1[38]), .B0(cout), .C0(n177_adj_5213), 
          .D0(d2[38]), .A1(d1[39]), .B1(cout), .C1(n174_adj_5212), .D1(d2[39]), 
          .CIN(n14939), .COUT(n14940), .S0(d2_71__N_490[38]), .S1(d2_71__N_490[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_3 (.A0(d1[36]), .B0(cout), .C0(n183_adj_5215), 
          .D0(d2[36]), .A1(d1[37]), .B1(cout), .C1(n180_adj_5214), .D1(d2[37]), 
          .CIN(n14938), .COUT(n14939), .S0(d2_71__N_490[36]), .S1(d2_71__N_490[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1517_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1517_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1517_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n14938));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1517_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1517_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1517_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1517_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_38 (.A0(d2_adj_5668[71]), .B0(d1_adj_5667[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14934), .S0(n78_adj_5562));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1568_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_36 (.A0(d2_adj_5668[69]), .B0(d1_adj_5667[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[70]), .B1(d1_adj_5667[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14933), .COUT(n14934), .S0(n84_adj_5564), 
          .S1(n81_adj_5563));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_34 (.A0(d2_adj_5668[67]), .B0(d1_adj_5667[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[68]), .B1(d1_adj_5667[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14932), .COUT(n14933), .S0(n90_adj_5566), 
          .S1(n87_adj_5565));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_32 (.A0(d2_adj_5668[65]), .B0(d1_adj_5667[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[66]), .B1(d1_adj_5667[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14931), .COUT(n14932), .S0(n96_adj_5568), 
          .S1(n93_adj_5567));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_30 (.A0(d2_adj_5668[63]), .B0(d1_adj_5667[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[64]), .B1(d1_adj_5667[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14930), .COUT(n14931), .S0(n102_adj_5570), 
          .S1(n99_adj_5569));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_28 (.A0(d2_adj_5668[61]), .B0(d1_adj_5667[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[62]), .B1(d1_adj_5667[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14929), .COUT(n14930), .S0(n108_adj_5572), 
          .S1(n105_adj_5571));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_26 (.A0(d2_adj_5668[59]), .B0(d1_adj_5667[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[60]), .B1(d1_adj_5667[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14928), .COUT(n14929), .S0(n114_adj_5574), 
          .S1(n111_adj_5573));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_24 (.A0(d2_adj_5668[57]), .B0(d1_adj_5667[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[58]), .B1(d1_adj_5667[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14927), .COUT(n14928), .S0(n120_adj_5576), 
          .S1(n117_adj_5575));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_22 (.A0(d2_adj_5668[55]), .B0(d1_adj_5667[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[56]), .B1(d1_adj_5667[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14926), .COUT(n14927), .S0(n126_adj_5578), 
          .S1(n123_adj_5577));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_20 (.A0(d2_adj_5668[53]), .B0(d1_adj_5667[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[54]), .B1(d1_adj_5667[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14925), .COUT(n14926), .S0(n132_adj_5580), 
          .S1(n129_adj_5579));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_18 (.A0(d2_adj_5668[51]), .B0(d1_adj_5667[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[52]), .B1(d1_adj_5667[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14924), .COUT(n14925), .S0(n138_adj_5582), 
          .S1(n135_adj_5581));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_16 (.A0(d2_adj_5668[49]), .B0(d1_adj_5667[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[50]), .B1(d1_adj_5667[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14923), .COUT(n14924), .S0(n144_adj_5584), 
          .S1(n141_adj_5583));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_14 (.A0(d2_adj_5668[47]), .B0(d1_adj_5667[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[48]), .B1(d1_adj_5667[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14922), .COUT(n14923), .S0(n150_adj_5586), 
          .S1(n147_adj_5585));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_12 (.A0(d2_adj_5668[45]), .B0(d1_adj_5667[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[46]), .B1(d1_adj_5667[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14921), .COUT(n14922), .S0(n156_adj_5588), 
          .S1(n153_adj_5587));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_10 (.A0(d2_adj_5668[43]), .B0(d1_adj_5667[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[44]), .B1(d1_adj_5667[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14920), .COUT(n14921), .S0(n162_adj_5590), 
          .S1(n159_adj_5589));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_8 (.A0(d2_adj_5668[41]), .B0(d1_adj_5667[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[42]), .B1(d1_adj_5667[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14919), .COUT(n14920), .S0(n168_adj_5592), 
          .S1(n165_adj_5591));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_6 (.A0(d2_adj_5668[39]), .B0(d1_adj_5667[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[40]), .B1(d1_adj_5667[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14918), .COUT(n14919), .S0(n174_adj_5594), 
          .S1(n171_adj_5593));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1568_add_4_4 (.A0(d2_adj_5668[37]), .B0(d1_adj_5667[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[38]), .B1(d1_adj_5667[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14917), .COUT(n14918), .S0(n180_adj_5596), 
          .S1(n177_adj_5595));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1568_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_4.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i2 (.D(n123_adj_5177), .CK(CIC1_out_clkSin), .Q(ISquare[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i2.GSR = "ENABLED";
    CCU2C _add_1_1568_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2_adj_5668[36]), .B1(d1_adj_5667[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14917), .S1(n183_adj_5597));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1568_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1568_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1568_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1568_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_38 (.A0(d_d9[35]), .B0(d9[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14916), .S1(cout_adj_5656));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1619_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_36 (.A0(d_d9[33]), .B0(d9[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[34]), .B1(d9[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14915), .COUT(n14916));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_34 (.A0(d_d9[31]), .B0(d9[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[32]), .B1(d9[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14914), .COUT(n14915));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_32 (.A0(d_d9[29]), .B0(d9[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[30]), .B1(d9[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14913), .COUT(n14914));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_30 (.A0(d_d9[27]), .B0(d9[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[28]), .B1(d9[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14912), .COUT(n14913));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_28 (.A0(d_d9[25]), .B0(d9[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[26]), .B1(d9[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14911), .COUT(n14912));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_26 (.A0(d_d9[23]), .B0(d9[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[24]), .B1(d9[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14910), .COUT(n14911));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_24 (.A0(d_d9[21]), .B0(d9[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[22]), .B1(d9[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14909), .COUT(n14910));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_22 (.A0(d_d9[19]), .B0(d9[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[20]), .B1(d9[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14908), .COUT(n14909));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_22.INJECT1_1 = "NO";
    LUT4 equal_298_i11_2_lut (.A(o_Rx_Byte[2]), .B(n17751), .Z(n11_adj_4566)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_298_i11_2_lut.init = 16'heeee;
    CCU2C _add_1_1619_add_4_14 (.A0(d_d9[11]), .B0(d9[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[12]), .B1(d9[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14904), .COUT(n14905));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_20 (.A0(d_d9[17]), .B0(d9[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[18]), .B1(d9[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14907), .COUT(n14908));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_10 (.A0(d_d9[7]), .B0(d9[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[8]), .B1(d9[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14902), .COUT(n14903));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_18 (.A0(d_d9[15]), .B0(d9[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[16]), .B1(d9[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14906), .COUT(n14907));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_8 (.A0(d_d9[5]), .B0(d9[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[6]), .B1(d9[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14901), .COUT(n14902));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_6 (.A0(d_d9[3]), .B0(d9[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[4]), .B1(d9[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14900), .COUT(n14901));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[0]), .B1(d9[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n14899));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1619_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_12 (.A0(d_d9[9]), .B0(d9[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[10]), .B1(d9[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14903), .COUT(n14904));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1619_add_4_16 (.A0(d_d9[13]), .B0(d9[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[14]), .B1(d9[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14905), .COUT(n14906));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_16.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i3 (.D(n120_adj_5176), .CK(CIC1_out_clkSin), .Q(ISquare[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i3.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i4 (.D(n117_adj_5175), .CK(CIC1_out_clkSin), .Q(ISquare[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i4.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i5 (.D(n114_adj_5174), .CK(CIC1_out_clkSin), .Q(ISquare[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i5.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i6 (.D(n111_adj_5173), .CK(CIC1_out_clkSin), .Q(ISquare[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i6.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i7 (.D(n108_adj_5172), .CK(CIC1_out_clkSin), .Q(ISquare[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i7.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i8 (.D(n105_adj_5171), .CK(CIC1_out_clkSin), .Q(ISquare[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i8.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i9 (.D(n102_adj_5170), .CK(CIC1_out_clkSin), .Q(ISquare[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i9.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i10 (.D(n99_adj_5169), .CK(CIC1_out_clkSin), .Q(ISquare[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i10.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i11 (.D(n96_adj_5168), .CK(CIC1_out_clkSin), .Q(ISquare[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i11.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i12 (.D(n93_adj_5167), .CK(CIC1_out_clkSin), .Q(ISquare[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i12.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i13 (.D(n90_adj_5166), .CK(CIC1_out_clkSin), .Q(ISquare[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i13.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i14 (.D(n87_adj_5165), .CK(CIC1_out_clkSin), .Q(ISquare[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i14.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i15 (.D(n84_adj_5164), .CK(CIC1_out_clkSin), .Q(ISquare[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i15.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i16 (.D(n81_adj_5163), .CK(CIC1_out_clkSin), .Q(ISquare[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i16.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i17 (.D(n78_adj_5162), .CK(CIC1_out_clkSin), .Q(ISquare[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i17.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i18 (.D(n75_adj_5161), .CK(CIC1_out_clkSin), .Q(ISquare[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i18.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i19 (.D(n72_adj_5160), .CK(CIC1_out_clkSin), .Q(ISquare[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i19.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i20 (.D(n69_adj_5159), .CK(CIC1_out_clkSin), .Q(ISquare[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i20.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i21 (.D(n66_adj_5158), .CK(CIC1_out_clkSin), .Q(ISquare[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i21.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i22 (.D(n63_adj_5157), .CK(CIC1_out_clkSin), .Q(ISquare[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i22.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i23 (.D(n60_adj_5156), .CK(CIC1_out_clkSin), .Q(ISquare[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i23.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i24 (.D(n57_adj_5155), .CK(CIC1_out_clkSin), .Q(ISquare[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i24.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i25 (.D(n54_adj_5154), .CK(CIC1_out_clkSin), .Q(ISquare[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_e3__i25.GSR = "ENABLED";
    CCU2C add_3645_45 (.A0(phase_inc_carrGen[42]), .B0(n13169), .C0(n2328), 
          .D0(n17621), .A1(phase_inc_carrGen[43]), .B1(n13169), .C1(n2327), 
          .D1(n3676), .CIN(n16354), .COUT(n16355), .S0(n197), .S1(n194));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_45.INIT0 = 16'h74b8;
    defparam add_3645_45.INIT1 = 16'h74b8;
    defparam add_3645_45.INJECT1_0 = "NO";
    defparam add_3645_45.INJECT1_1 = "NO";
    CCU2C add_3645_43 (.A0(phase_inc_carrGen[40]), .B0(n13169), .C0(n2330), 
          .D0(n3656), .A1(phase_inc_carrGen[41]), .B1(n13169), .C1(n12140), 
          .D1(n3676), .CIN(n16353), .COUT(n16354), .S0(n203), .S1(n200));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_43.INIT0 = 16'h74b8;
    defparam add_3645_43.INIT1 = 16'h74b8;
    defparam add_3645_43.INJECT1_0 = "NO";
    defparam add_3645_43.INJECT1_1 = "NO";
    CCU2C add_3645_41 (.A0(phase_inc_carrGen[38]), .B0(n13169), .C0(n2332), 
          .D0(n3659), .A1(phase_inc_carrGen[39]), .B1(n13169), .C1(n2331), 
          .D1(n3659), .CIN(n16352), .COUT(n16353), .S0(n209_adj_4997), 
          .S1(n206));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_41.INIT0 = 16'h74b8;
    defparam add_3645_41.INIT1 = 16'h74b8;
    defparam add_3645_41.INJECT1_0 = "NO";
    defparam add_3645_41.INJECT1_1 = "NO";
    CCU2C add_3645_39 (.A0(phase_inc_carrGen[36]), .B0(n13169), .C0(n2334), 
          .D0(n17622), .A1(phase_inc_carrGen[37]), .B1(n13169), .C1(n2333), 
          .D1(n3677), .CIN(n16351), .COUT(n16352), .S0(n215), .S1(n212));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_39.INIT0 = 16'h74b8;
    defparam add_3645_39.INIT1 = 16'h74b8;
    defparam add_3645_39.INJECT1_0 = "NO";
    defparam add_3645_39.INJECT1_1 = "NO";
    CCU2C add_3645_37 (.A0(phase_inc_carrGen[34]), .B0(n13169), .C0(n2336), 
          .D0(n17622), .A1(phase_inc_carrGen[35]), .B1(n13169), .C1(n2335), 
          .D1(n3659), .CIN(n16350), .COUT(n16351), .S0(n221), .S1(n218));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_37.INIT0 = 16'h74b8;
    defparam add_3645_37.INIT1 = 16'h74b8;
    defparam add_3645_37.INJECT1_0 = "NO";
    defparam add_3645_37.INJECT1_1 = "NO";
    CCU2C add_3645_35 (.A0(phase_inc_carrGen[32]), .B0(n13169), .C0(n2338), 
          .D0(n3656), .A1(phase_inc_carrGen[33]), .B1(n13169), .C1(n2337), 
          .D1(n3677), .CIN(n16349), .COUT(n16350), .S0(n227), .S1(n224));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_35.INIT0 = 16'h74b8;
    defparam add_3645_35.INIT1 = 16'h74b8;
    defparam add_3645_35.INJECT1_0 = "NO";
    defparam add_3645_35.INJECT1_1 = "NO";
    CCU2C add_3645_33 (.A0(phase_inc_carrGen[30]), .B0(n13169), .C0(n2340), 
          .D0(n3656), .A1(phase_inc_carrGen[31]), .B1(n13169), .C1(n2339), 
          .D1(n3691), .CIN(n16348), .COUT(n16349), .S0(n233), .S1(n230));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_33.INIT0 = 16'h74b8;
    defparam add_3645_33.INIT1 = 16'h74b8;
    defparam add_3645_33.INJECT1_0 = "NO";
    defparam add_3645_33.INJECT1_1 = "NO";
    CCU2C add_3645_31 (.A0(phase_inc_carrGen[28]), .B0(n13169), .C0(n2342), 
          .D0(n3676), .A1(phase_inc_carrGen[29]), .B1(n13169), .C1(n2341), 
          .D1(n17621), .CIN(n16347), .COUT(n16348), .S0(n239), .S1(n236));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_31.INIT0 = 16'h74b8;
    defparam add_3645_31.INIT1 = 16'h74b8;
    defparam add_3645_31.INJECT1_0 = "NO";
    defparam add_3645_31.INJECT1_1 = "NO";
    CCU2C add_3645_29 (.A0(phase_inc_carrGen[26]), .B0(n13169), .C0(n2344), 
          .D0(n3659), .A1(phase_inc_carrGen[27]), .B1(n13169), .C1(n2343), 
          .D1(n3677), .CIN(n16346), .COUT(n16347), .S0(n245), .S1(n242));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_29.INIT0 = 16'h74b8;
    defparam add_3645_29.INIT1 = 16'h74b8;
    defparam add_3645_29.INJECT1_0 = "NO";
    defparam add_3645_29.INJECT1_1 = "NO";
    CCU2C add_3645_27 (.A0(phase_inc_carrGen[24]), .B0(n13169), .C0(n2346), 
          .D0(n3659), .A1(phase_inc_carrGen[25]), .B1(n13169), .C1(n2345), 
          .D1(n3659), .CIN(n16345), .COUT(n16346), .S0(n251), .S1(n248));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_27.INIT0 = 16'h74b8;
    defparam add_3645_27.INIT1 = 16'h74b8;
    defparam add_3645_27.INJECT1_0 = "NO";
    defparam add_3645_27.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15611), .S1(MixerOutSin_11__N_236[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(41[26:33])
    defparam _add_1_1454_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1454_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1454_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_1.INJECT1_1 = "NO";
    CCU2C add_3645_25 (.A0(phase_inc_carrGen[22]), .B0(n13169), .C0(n2348), 
          .D0(n17622), .A1(phase_inc_carrGen[23]), .B1(n13169), .C1(n2347), 
          .D1(n17621), .CIN(n16344), .COUT(n16345), .S0(n257), .S1(n254));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_25.INIT0 = 16'h74b8;
    defparam add_3645_25.INIT1 = 16'h74b8;
    defparam add_3645_25.INJECT1_0 = "NO";
    defparam add_3645_25.INJECT1_1 = "NO";
    CCU2C add_3645_23 (.A0(phase_inc_carrGen[20]), .B0(n13169), .C0(n2350), 
          .D0(n3659), .A1(phase_inc_carrGen[21]), .B1(n13169), .C1(n2349), 
          .D1(n3656), .CIN(n16343), .COUT(n16344), .S0(n263), .S1(n260));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_23.INIT0 = 16'h74b8;
    defparam add_3645_23.INIT1 = 16'h74b8;
    defparam add_3645_23.INJECT1_0 = "NO";
    defparam add_3645_23.INJECT1_1 = "NO";
    CCU2C add_3645_21 (.A0(phase_inc_carrGen[18]), .B0(n13169), .C0(n2352), 
          .D0(n17621), .A1(phase_inc_carrGen[19]), .B1(n13169), .C1(n12138), 
          .D1(n3677), .CIN(n16342), .COUT(n16343), .S0(n269), .S1(n266));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_21.INIT0 = 16'h74b8;
    defparam add_3645_21.INIT1 = 16'h74b8;
    defparam add_3645_21.INJECT1_0 = "NO";
    defparam add_3645_21.INJECT1_1 = "NO";
    CCU2C add_3645_19 (.A0(phase_inc_carrGen[16]), .B0(n13169), .C0(n2354), 
          .D0(n3691), .A1(phase_inc_carrGen[17]), .B1(n13169), .C1(n12136), 
          .D1(n11690), .CIN(n16341), .COUT(n16342), .S0(n275), .S1(n272));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_19.INIT0 = 16'h74b8;
    defparam add_3645_19.INIT1 = 16'h74b8;
    defparam add_3645_19.INJECT1_0 = "NO";
    defparam add_3645_19.INJECT1_1 = "NO";
    CCU2C add_3645_17 (.A0(phase_inc_carrGen[14]), .B0(n13169), .C0(n2356), 
          .D0(n17622), .A1(phase_inc_carrGen[15]), .B1(n13169), .C1(n2355), 
          .D1(n3677), .CIN(n16340), .COUT(n16341), .S0(n281), .S1(n278));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_17.INIT0 = 16'h74b8;
    defparam add_3645_17.INIT1 = 16'h74b8;
    defparam add_3645_17.INJECT1_0 = "NO";
    defparam add_3645_17.INJECT1_1 = "NO";
    CCU2C add_3645_15 (.A0(phase_inc_carrGen[12]), .B0(n13169), .C0(n2358), 
          .D0(n17622), .A1(phase_inc_carrGen[13]), .B1(n13169), .C1(n12134), 
          .D1(n3691), .CIN(n16339), .COUT(n16340), .S0(n287), .S1(n284));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_15.INIT0 = 16'h74b8;
    defparam add_3645_15.INIT1 = 16'h74b8;
    defparam add_3645_15.INJECT1_0 = "NO";
    defparam add_3645_15.INJECT1_1 = "NO";
    CCU2C add_3645_13 (.A0(phase_inc_carrGen[10]), .B0(n13169), .C0(n2360), 
          .D0(n3691), .A1(phase_inc_carrGen[11]), .B1(n13169), .C1(n2359), 
          .D1(n3659), .CIN(n16338), .COUT(n16339), .S0(n293), .S1(n290));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_13.INIT0 = 16'h74b8;
    defparam add_3645_13.INIT1 = 16'h74b8;
    defparam add_3645_13.INJECT1_0 = "NO";
    defparam add_3645_13.INJECT1_1 = "NO";
    CCU2C add_3645_11 (.A0(phase_inc_carrGen[8]), .B0(n13169), .C0(n2362), 
          .D0(n3676), .A1(phase_inc_carrGen[9]), .B1(n13169), .C1(n2361), 
          .D1(n17621), .CIN(n16337), .COUT(n16338), .S0(n299), .S1(n296));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_11.INIT0 = 16'h74b8;
    defparam add_3645_11.INIT1 = 16'h74b8;
    defparam add_3645_11.INJECT1_0 = "NO";
    defparam add_3645_11.INJECT1_1 = "NO";
    CCU2C add_3645_9 (.A0(phase_inc_carrGen[6]), .B0(n13169), .C0(n12132), 
          .D0(n3677), .A1(phase_inc_carrGen[7]), .B1(n13169), .C1(n2363), 
          .D1(n17621), .CIN(n16336), .COUT(n16337), .S0(n305), .S1(n302));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_9.INIT0 = 16'h74b8;
    defparam add_3645_9.INIT1 = 16'h74b8;
    defparam add_3645_9.INJECT1_0 = "NO";
    defparam add_3645_9.INJECT1_1 = "NO";
    CCU2C add_3645_7 (.A0(phase_inc_carrGen[4]), .B0(n13169), .C0(n2366), 
          .D0(n3677), .A1(phase_inc_carrGen[5]), .B1(n13169), .C1(n2365), 
          .D1(n3677), .CIN(n16335), .COUT(n16336), .S0(n311), .S1(n308));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_7.INIT0 = 16'h74b8;
    defparam add_3645_7.INIT1 = 16'h74b8;
    defparam add_3645_7.INJECT1_0 = "NO";
    defparam add_3645_7.INJECT1_1 = "NO";
    CCU2C add_3645_5 (.A0(phase_inc_carrGen[2]), .B0(n13169), .C0(n2368), 
          .D0(n11690), .A1(phase_inc_carrGen[3]), .B1(n13169), .C1(n2367), 
          .D1(n11690), .CIN(n16334), .COUT(n16335), .S0(n317), .S1(n314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_5.INIT0 = 16'h74b8;
    defparam add_3645_5.INIT1 = 16'h74b8;
    defparam add_3645_5.INJECT1_0 = "NO";
    defparam add_3645_5.INJECT1_1 = "NO";
    CCU2C add_3645_3 (.A0(phase_inc_carrGen[0]), .B0(n13169), .C0(n2636), 
          .D0(n17621), .A1(phase_inc_carrGen[1]), .B1(n13169), .C1(n2369), 
          .D1(n3691), .CIN(n16333), .COUT(n16334), .S0(n323), .S1(n320));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_3.INIT0 = 16'h74b8;
    defparam add_3645_3.INIT1 = 16'h74b8;
    defparam add_3645_3.INJECT1_0 = "NO";
    defparam add_3645_3.INJECT1_1 = "NO";
    CCU2C add_3645_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n17618), .B1(n12966), .C1(o_Rx_Byte[4]), .D1(n2823), .COUT(n16333));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam add_3645_1.INIT0 = 16'h0000;
    defparam add_3645_1.INIT1 = 16'hf7ff;
    defparam add_3645_1.INJECT1_0 = "NO";
    defparam add_3645_1.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_38 (.A0(d5[71]), .B0(d4[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15610), .S0(n78_adj_5384));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1562_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_38.INJECT1_1 = "NO";
    CCU2C add_3646_17 (.A0(d_out_d_11__N_1877), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1877), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16328), .S0(n51_adj_5255), 
          .S1(d_out_d_11__N_1880[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_17.INIT0 = 16'h666a;
    defparam add_3646_17.INIT1 = 16'h666a;
    defparam add_3646_17.INJECT1_0 = "NO";
    defparam add_3646_17.INJECT1_1 = "NO";
    CCU2C add_3646_15 (.A0(d_out_d_11__N_1878[17]), .B0(n55), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n52), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16327), .COUT(n16328), .S0(n57_adj_5257), 
          .S1(n54_adj_5256));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_15.INIT0 = 16'h9995;
    defparam add_3646_15.INIT1 = 16'h9995;
    defparam add_3646_15.INJECT1_0 = "NO";
    defparam add_3646_15.INJECT1_1 = "NO";
    CCU2C add_3646_13 (.A0(d_out_d_11__N_1878[17]), .B0(n61), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n58), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16326), .COUT(n16327), .S0(n63_adj_5259), 
          .S1(n60_adj_5258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_13.INIT0 = 16'h9995;
    defparam add_3646_13.INIT1 = 16'h9995;
    defparam add_3646_13.INJECT1_0 = "NO";
    defparam add_3646_13.INJECT1_1 = "NO";
    CCU2C add_3646_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1878[17]), .C0(n67_adj_5379), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n64_adj_5378), .D1(VCC_net), .CIN(n16325), .COUT(n16326), 
          .S0(n69_adj_5261), .S1(n66_adj_5260));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_11.INIT0 = 16'h6969;
    defparam add_3646_11.INIT1 = 16'h6969;
    defparam add_3646_11.INJECT1_0 = "NO";
    defparam add_3646_11.INJECT1_1 = "NO";
    CCU2C add_3646_9 (.A0(d_out_d_11__N_1878[17]), .B0(n73), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n70), .D1(VCC_net), .CIN(n16324), .COUT(n16325), .S0(n75_adj_5263), 
          .S1(n72_adj_5262));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_9.INIT0 = 16'h9995;
    defparam add_3646_9.INIT1 = 16'h6969;
    defparam add_3646_9.INJECT1_0 = "NO";
    defparam add_3646_9.INJECT1_1 = "NO";
    CCU2C add_3646_7 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1878[17]), 
          .C0(n79_adj_5381), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(n17635), .C1(n76_adj_5380), .D1(VCC_net), .CIN(n16323), 
          .COUT(n16324), .S0(n81_adj_5265), .S1(n78_adj_5264));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_7.INIT0 = 16'h9696;
    defparam add_3646_7.INIT1 = 16'h6969;
    defparam add_3646_7.INJECT1_0 = "NO";
    defparam add_3646_7.INJECT1_1 = "NO";
    CCU2C add_3646_5 (.A0(n85_adj_5383), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1878[17]), .C1(n82_adj_5382), 
          .D1(VCC_net), .CIN(n16322), .COUT(n16323), .S0(n87_adj_5267), 
          .S1(n84_adj_5266));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_5.INIT0 = 16'haaa0;
    defparam add_3646_5.INIT1 = 16'h9696;
    defparam add_3646_5.INJECT1_0 = "NO";
    defparam add_3646_5.INJECT1_1 = "NO";
    CCU2C add_3646_3 (.A0(d_out_d_11__N_1878[17]), .B0(ISquare[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16321), .COUT(n16322), .S1(n90_adj_5268));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_3.INIT0 = 16'h666a;
    defparam add_3646_3.INIT1 = 16'h555f;
    defparam add_3646_3.INJECT1_0 = "NO";
    defparam add_3646_3.INJECT1_1 = "NO";
    CCU2C add_3646_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16321));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3646_1.INIT0 = 16'h0000;
    defparam add_3646_1.INIT1 = 16'haaaf;
    defparam add_3646_1.INJECT1_0 = "NO";
    defparam add_3646_1.INJECT1_1 = "NO";
    CCU2C add_3641_19 (.A0(d_out_d_11__N_1884[17]), .B0(n48_adj_5474), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n45_adj_5473), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16315), .S0(n45_adj_5421), 
          .S1(d_out_d_11__N_1886[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_19.INIT0 = 16'h9995;
    defparam add_3641_19.INIT1 = 16'h9995;
    defparam add_3641_19.INJECT1_0 = "NO";
    defparam add_3641_19.INJECT1_1 = "NO";
    CCU2C add_3641_17 (.A0(d_out_d_11__N_1884[17]), .B0(n54_adj_5476), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n51_adj_5475), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16314), .COUT(n16315), .S0(n51_adj_5423), 
          .S1(n48_adj_5422));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_17.INIT0 = 16'h9995;
    defparam add_3641_17.INIT1 = 16'h9995;
    defparam add_3641_17.INJECT1_0 = "NO";
    defparam add_3641_17.INJECT1_1 = "NO";
    CCU2C add_3641_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n60_adj_5478), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n57_adj_5477), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16313), .COUT(n16314), .S0(n57_adj_5425), 
          .S1(n54_adj_5424));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_15.INIT0 = 16'h6969;
    defparam add_3641_15.INIT1 = 16'h9995;
    defparam add_3641_15.INJECT1_0 = "NO";
    defparam add_3641_15.INJECT1_1 = "NO";
    CCU2C add_3641_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n66_adj_5480), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1884[17]), 
          .C1(n63_adj_5479), .D1(VCC_net), .CIN(n16312), .COUT(n16313), 
          .S0(n63_adj_5427), .S1(n60_adj_5426));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_13.INIT0 = 16'h6969;
    defparam add_3641_13.INIT1 = 16'h6969;
    defparam add_3641_13.INJECT1_0 = "NO";
    defparam add_3641_13.INJECT1_1 = "NO";
    CCU2C add_3641_11 (.A0(d_out_d_11__N_1884[17]), .B0(n17635), .C0(n72_adj_5482), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n69_adj_5481), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16311), .COUT(n16312), .S0(n69_adj_5429), 
          .S1(n66_adj_5428));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_11.INIT0 = 16'h6969;
    defparam add_3641_11.INIT1 = 16'h9995;
    defparam add_3641_11.INJECT1_0 = "NO";
    defparam add_3641_11.INJECT1_1 = "NO";
    CCU2C add_3641_9 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n78_adj_5484), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n75_adj_5483), .D1(VCC_net), 
          .CIN(n16310), .COUT(n16311), .S0(n75_adj_5431), .S1(n72_adj_5430));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_9.INIT0 = 16'h9696;
    defparam add_3641_9.INIT1 = 16'h9696;
    defparam add_3641_9.INJECT1_0 = "NO";
    defparam add_3641_9.INJECT1_1 = "NO";
    CCU2C add_3641_7 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n84_adj_5486), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n81_adj_5485), .D1(VCC_net), 
          .CIN(n16309), .COUT(n16310), .S0(n81_adj_5433), .S1(n78_adj_5432));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_7.INIT0 = 16'h9696;
    defparam add_3641_7.INIT1 = 16'h9696;
    defparam add_3641_7.INJECT1_0 = "NO";
    defparam add_3641_7.INJECT1_1 = "NO";
    CCU2C add_3641_5 (.A0(n90_adj_5488), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(d_out_d_11__N_1884[17]), .C1(n87_adj_5487), 
          .D1(VCC_net), .CIN(n16308), .COUT(n16309), .S0(n87_adj_5435), 
          .S1(n84_adj_5434));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_5.INIT0 = 16'haaa0;
    defparam add_3641_5.INIT1 = 16'h9696;
    defparam add_3641_5.INJECT1_0 = "NO";
    defparam add_3641_5.INJECT1_1 = "NO";
    CCU2C add_3641_3 (.A0(d_out_d_11__N_1884[17]), .B0(ISquare[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16307), .COUT(n16308), .S1(n90_adj_5436));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_3.INIT0 = 16'h666a;
    defparam add_3641_3.INIT1 = 16'h555f;
    defparam add_3641_3.INJECT1_0 = "NO";
    defparam add_3641_3.INJECT1_1 = "NO";
    CCU2C add_3641_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16307));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3641_1.INIT0 = 16'h0000;
    defparam add_3641_1.INIT1 = 16'haaaf;
    defparam add_3641_1.INJECT1_0 = "NO";
    defparam add_3641_1.INJECT1_1 = "NO";
    CCU2C add_3642_13 (.A0(d_out_d_11__N_1873), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1873), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16301), .S0(n48_adj_5552), 
          .S1(d_out_d_11__N_1876[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_13.INIT0 = 16'h666a;
    defparam add_3642_13.INIT1 = 16'h666a;
    defparam add_3642_13.INJECT1_0 = "NO";
    defparam add_3642_13.INJECT1_1 = "NO";
    CCU2C add_3642_11 (.A0(d_out_d_11__N_1874[17]), .B0(n47), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n44), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16300), .COUT(n16301), .S0(n54_adj_5554), 
          .S1(n51_adj_5553));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_11.INIT0 = 16'h9995;
    defparam add_3642_11.INIT1 = 16'h9995;
    defparam add_3642_11.INJECT1_0 = "NO";
    defparam add_3642_11.INJECT1_1 = "NO";
    CCU2C add_3642_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1874[17]), .C0(n53), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n50), .D1(VCC_net), .CIN(n16299), .COUT(n16300), .S0(n60_adj_5556), 
          .S1(n57_adj_5555));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_9.INIT0 = 16'h6969;
    defparam add_3642_9.INIT1 = 16'h6969;
    defparam add_3642_9.INJECT1_0 = "NO";
    defparam add_3642_9.INJECT1_1 = "NO";
    CCU2C add_3642_7 (.A0(d_out_d_11__N_1874[17]), .B0(n59), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n56), .D1(VCC_net), .CIN(n16298), .COUT(n16299), .S0(n66_adj_5558), 
          .S1(n63_adj_5557));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_7.INIT0 = 16'h9995;
    defparam add_3642_7.INIT1 = 16'h6969;
    defparam add_3642_7.INJECT1_0 = "NO";
    defparam add_3642_7.INJECT1_1 = "NO";
    CCU2C add_3642_5 (.A0(n65), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(n17635), .C1(n62), .D1(VCC_net), 
          .CIN(n16297), .COUT(n16298), .S0(n72_adj_5560), .S1(n69_adj_5559));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_5.INIT0 = 16'haaa0;
    defparam add_3642_5.INIT1 = 16'h6969;
    defparam add_3642_5.INJECT1_0 = "NO";
    defparam add_3642_5.INJECT1_1 = "NO";
    CCU2C add_3642_3 (.A0(d_out_d_11__N_1874[17]), .B0(ISquare[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16296), .COUT(n16297), .S1(n75_adj_5561));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_3.INIT0 = 16'h666a;
    defparam add_3642_3.INIT1 = 16'h555f;
    defparam add_3642_3.INJECT1_0 = "NO";
    defparam add_3642_3.INJECT1_1 = "NO";
    CCU2C add_3642_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16296));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3642_1.INIT0 = 16'h0000;
    defparam add_3642_1.INIT1 = 16'haaaf;
    defparam add_3642_1.INJECT1_0 = "NO";
    defparam add_3642_1.INJECT1_1 = "NO";
    CCU2C add_3635_19 (.A0(d_out_d_11__N_1888[17]), .B0(n48_adj_5537), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n45_adj_5536), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16290), .S0(n45_adj_5505), 
          .S1(d_out_d_11__N_1890[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_19.INIT0 = 16'h9995;
    defparam add_3635_19.INIT1 = 16'h9995;
    defparam add_3635_19.INJECT1_0 = "NO";
    defparam add_3635_19.INJECT1_1 = "NO";
    CCU2C add_3635_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n54_adj_5539), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n51_adj_5538), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16289), .COUT(n16290), .S0(n51_adj_5507), 
          .S1(n48_adj_5506));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_17.INIT0 = 16'h6969;
    defparam add_3635_17.INIT1 = 16'h9995;
    defparam add_3635_17.INJECT1_0 = "NO";
    defparam add_3635_17.INJECT1_1 = "NO";
    CCU2C add_3635_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n60_adj_5541), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1888[17]), 
          .C1(n57_adj_5540), .D1(VCC_net), .CIN(n16288), .COUT(n16289), 
          .S0(n57_adj_5509), .S1(n54_adj_5508));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_15.INIT0 = 16'h6969;
    defparam add_3635_15.INIT1 = 16'h6969;
    defparam add_3635_15.INJECT1_0 = "NO";
    defparam add_3635_15.INJECT1_1 = "NO";
    CCU2C add_3635_13 (.A0(d_out_d_11__N_1888[17]), .B0(n17635), .C0(n66_adj_5543), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n63_adj_5542), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16287), .COUT(n16288), .S0(n63_adj_5511), 
          .S1(n60_adj_5510));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_13.INIT0 = 16'h6969;
    defparam add_3635_13.INIT1 = 16'h9995;
    defparam add_3635_13.INJECT1_0 = "NO";
    defparam add_3635_13.INJECT1_1 = "NO";
    CCU2C add_3635_11 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n72_adj_5545), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n69_adj_5544), .D1(VCC_net), 
          .CIN(n16286), .COUT(n16287), .S0(n69_adj_5513), .S1(n66_adj_5512));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_11.INIT0 = 16'h9696;
    defparam add_3635_11.INIT1 = 16'h9696;
    defparam add_3635_11.INJECT1_0 = "NO";
    defparam add_3635_11.INJECT1_1 = "NO";
    CCU2C add_3635_9 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n78_adj_5547), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n75_adj_5546), .D1(VCC_net), 
          .CIN(n16285), .COUT(n16286), .S0(n75_adj_5515), .S1(n72_adj_5514));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_9.INIT0 = 16'h9696;
    defparam add_3635_9.INIT1 = 16'h9696;
    defparam add_3635_9.INJECT1_0 = "NO";
    defparam add_3635_9.INJECT1_1 = "NO";
    CCU2C add_3635_7 (.A0(d_out_d_11__N_1884[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n84_adj_5549), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n81_adj_5548), .D1(VCC_net), 
          .CIN(n16284), .COUT(n16285), .S0(n81_adj_5517), .S1(n78_adj_5516));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_7.INIT0 = 16'h9696;
    defparam add_3635_7.INIT1 = 16'h9696;
    defparam add_3635_7.INJECT1_0 = "NO";
    defparam add_3635_7.INJECT1_1 = "NO";
    CCU2C add_3635_5 (.A0(n90_adj_5551), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(d_out_d_11__N_1888[17]), .C1(n87_adj_5550), 
          .D1(VCC_net), .CIN(n16283), .COUT(n16284), .S0(n87_adj_5519), 
          .S1(n84_adj_5518));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_5.INIT0 = 16'haaa0;
    defparam add_3635_5.INIT1 = 16'h9696;
    defparam add_3635_5.INJECT1_0 = "NO";
    defparam add_3635_5.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_8 (.A0(d_d7_adj_5675[41]), .B0(d7_adj_5674[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[42]), .B1(d7_adj_5674[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16137), .COUT(n16138), .S0(n168_adj_5335), 
          .S1(n165_adj_5334));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_8.INJECT1_1 = "NO";
    CCU2C add_3635_3 (.A0(d_out_d_11__N_1888[17]), .B0(ISquare[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16282), .COUT(n16283), .S1(n90_adj_5520));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_3.INIT0 = 16'h666a;
    defparam add_3635_3.INIT1 = 16'h555f;
    defparam add_3635_3.INJECT1_0 = "NO";
    defparam add_3635_3.INJECT1_1 = "NO";
    CCU2C add_3635_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3635_1.INIT0 = 16'h0000;
    defparam add_3635_1.INIT1 = 16'haaaf;
    defparam add_3635_1.INJECT1_0 = "NO";
    defparam add_3635_1.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_6 (.A0(d_d7_adj_5675[39]), .B0(d7_adj_5674[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[40]), .B1(d7_adj_5674[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16136), .COUT(n16137), .S0(n174_adj_5337), 
          .S1(n171_adj_5336));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_6.INJECT1_1 = "NO";
    CCU2C add_3643_11 (.A0(ISquare[31]), .B0(n17642), .C0(n17635), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n17642), .C1(n17635), .D1(VCC_net), 
          .CIN(n16276), .S0(n44), .S1(d_out_d_11__N_1874[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3643_11.INIT0 = 16'he1e1;
    defparam add_3643_11.INIT1 = 16'he1e1;
    defparam add_3643_11.INJECT1_0 = "NO";
    defparam add_3643_11.INJECT1_1 = "NO";
    CCU2C add_3643_9 (.A0(n17635), .B0(ISquare[31]), .C0(ISquare[23]), 
          .D0(ISquare[22]), .A1(n40), .B1(n14874), .C1(n209), .D1(ISquare[31]), 
          .CIN(n16275), .COUT(n16276), .S0(n50), .S1(n47));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3643_9.INIT0 = 16'h6665;
    defparam add_3643_9.INIT1 = 16'h556a;
    defparam add_3643_9.INJECT1_0 = "NO";
    defparam add_3643_9.INJECT1_1 = "NO";
    CCU2C add_3643_7 (.A0(n49), .B0(ISquare[31]), .C0(ISquare[23]), .D0(ISquare[22]), 
          .A1(n17642), .B1(ISquare[31]), .C1(ISquare[23]), .D1(ISquare[22]), 
          .CIN(n16274), .COUT(n16275), .S0(n56), .S1(n53));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3643_7.INIT0 = 16'h999a;
    defparam add_3643_7.INIT1 = 16'haaa9;
    defparam add_3643_7.INJECT1_0 = "NO";
    defparam add_3643_7.INJECT1_1 = "NO";
    CCU2C add_3643_5 (.A0(ISquare[22]), .B0(ISquare[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[23]), .B1(ISquare[22]), .C1(ISquare[31]), 
          .D1(n14874), .CIN(n16273), .COUT(n16274), .S0(n62), .S1(n59));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3643_5.INIT0 = 16'h9999;
    defparam add_3643_5.INIT1 = 16'heee1;
    defparam add_3643_5.INJECT1_0 = "NO";
    defparam add_3643_5.INJECT1_1 = "NO";
    CCU2C add_3643_3 (.A0(ISquare[31]), .B0(n17642), .C0(ISquare[20]), 
          .D0(VCC_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16272), .COUT(n16273), .S1(n65));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3643_3.INIT0 = 16'he1e1;
    defparam add_3643_3.INIT1 = 16'h555f;
    defparam add_3643_3.INJECT1_0 = "NO";
    defparam add_3643_3.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_4 (.A0(d_d7_adj_5675[37]), .B0(d7_adj_5674[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5675[38]), .B1(d7_adj_5674[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16135), .COUT(n16136), .S0(n180_adj_5339), 
          .S1(n177_adj_5338));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1628_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_4.INJECT1_1 = "NO";
    CCU2C add_3643_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[22]), .B1(ISquare[23]), .C1(n209), .D1(ISquare[31]), 
          .COUT(n16272));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3643_1.INIT0 = 16'h0000;
    defparam add_3643_1.INIT1 = 16'h001f;
    defparam add_3643_1.INJECT1_0 = "NO";
    defparam add_3643_1.INJECT1_1 = "NO";
    CCU2C add_3638_19 (.A0(d_out_d_11__N_1890[17]), .B0(n48_adj_5506), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n45_adj_5505), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16266), .S0(n912), .S1(d_out_d_11__N_1892[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_19.INIT0 = 16'h9995;
    defparam add_3638_19.INIT1 = 16'h9995;
    defparam add_3638_19.INJECT1_0 = "NO";
    defparam add_3638_19.INJECT1_1 = "NO";
    CCU2C add_3638_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1890[17]), .C0(n54_adj_5508), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n51_adj_5507), .D1(VCC_net), .CIN(n16265), .COUT(n16266), 
          .S0(n914), .S1(n913));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_17.INIT0 = 16'h6969;
    defparam add_3638_17.INIT1 = 16'h6969;
    defparam add_3638_17.INJECT1_0 = "NO";
    defparam add_3638_17.INJECT1_1 = "NO";
    CCU2C add_3638_15 (.A0(d_out_d_11__N_1890[17]), .B0(n60_adj_5510), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n57_adj_5509), .D1(VCC_net), .CIN(n16264), .COUT(n16265), 
          .S0(n916), .S1(n915));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_15.INIT0 = 16'h9995;
    defparam add_3638_15.INIT1 = 16'h6969;
    defparam add_3638_15.INJECT1_0 = "NO";
    defparam add_3638_15.INJECT1_1 = "NO";
    CCU2C add_3638_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n66_adj_5512), .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), 
          .B1(n17635), .C1(n63_adj_5511), .D1(VCC_net), .CIN(n16263), 
          .COUT(n16264), .S0(n918), .S1(n917));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_13.INIT0 = 16'h9696;
    defparam add_3638_13.INIT1 = 16'h6969;
    defparam add_3638_13.INJECT1_0 = "NO";
    defparam add_3638_13.INJECT1_1 = "NO";
    CCU2C add_3638_11 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n72_adj_5514), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n69_adj_5513), .D1(VCC_net), 
          .CIN(n16262), .COUT(n16263), .S0(n920), .S1(n919));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_11.INIT0 = 16'h9696;
    defparam add_3638_11.INIT1 = 16'h9696;
    defparam add_3638_11.INJECT1_0 = "NO";
    defparam add_3638_11.INJECT1_1 = "NO";
    CCU2C _add_1_1628_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5675[36]), .B1(d7_adj_5674[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16135), .S1(n183_adj_5340));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1628_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1628_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1628_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1628_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_38 (.A0(d_d6[35]), .B0(d6[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16134), .S0(d7_71__N_1531[35]), .S1(cout_adj_5341));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1523_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_36 (.A0(d_d6[33]), .B0(d6[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[34]), .B1(d6[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16133), .COUT(n16134), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_34 (.A0(d_d6[31]), .B0(d6[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[32]), .B1(d6[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16132), .COUT(n16133), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_32 (.A0(d_d6[29]), .B0(d6[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[30]), .B1(d6[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16131), .COUT(n16132), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_30 (.A0(d_d6[27]), .B0(d6[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[28]), .B1(d6[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16130), .COUT(n16131), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_28 (.A0(d_d6[25]), .B0(d6[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[26]), .B1(d6[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16129), .COUT(n16130), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_26 (.A0(d_d6[23]), .B0(d6[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[24]), .B1(d6[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16128), .COUT(n16129), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_24 (.A0(d_d6[21]), .B0(d6[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[22]), .B1(d6[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16127), .COUT(n16128), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_22 (.A0(d_d6[19]), .B0(d6[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[20]), .B1(d6[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16126), .COUT(n16127), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_20 (.A0(d_d6[17]), .B0(d6[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[18]), .B1(d6[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16125), .COUT(n16126), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_18 (.A0(d_d6[15]), .B0(d6[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[16]), .B1(d6[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16124), .COUT(n16125), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_16 (.A0(d_d6[13]), .B0(d6[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[14]), .B1(d6[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16123), .COUT(n16124), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_14 (.A0(d_d6[11]), .B0(d6[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[12]), .B1(d6[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16122), .COUT(n16123), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_12 (.A0(d_d6[9]), .B0(d6[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[10]), .B1(d6[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16121), .COUT(n16122), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_10 (.A0(d_d6[7]), .B0(d6[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[8]), .B1(d6[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16120), .COUT(n16121), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_8 (.A0(d_d6[5]), .B0(d6[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[6]), .B1(d6[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16119), .COUT(n16120), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_6 (.A0(d_d6[3]), .B0(d6[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[4]), .B1(d6[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16118), .COUT(n16119), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_4 (.A0(d_d6[1]), .B0(d6[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[2]), .B1(d6[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16117), .COUT(n16118), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1523_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1523_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[0]), .B1(d6[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16117), .S1(d7_71__N_1531[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1523_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1523_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1523_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1523_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_37 (.A0(d_tmp[70]), .B0(cout_adj_5217), .C0(n81_adj_4962), 
          .D0(n3_adj_4763), .A1(d_tmp[71]), .B1(cout_adj_5217), .C1(n78_adj_4961), 
          .D1(n2_adj_4764), .CIN(n16115), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_35 (.A0(d_tmp[68]), .B0(cout_adj_5217), .C0(n87_adj_4964), 
          .D0(n5_adj_4761), .A1(d_tmp[69]), .B1(cout_adj_5217), .C1(n84_adj_4963), 
          .D1(n4_adj_4762), .CIN(n16114), .COUT(n16115), .S0(d6_71__N_1459[68]), 
          .S1(d6_71__N_1459[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_33 (.A0(d_tmp[66]), .B0(cout_adj_5217), .C0(n93_adj_4966), 
          .D0(n7_adj_4759), .A1(d_tmp[67]), .B1(cout_adj_5217), .C1(n90_adj_4965), 
          .D1(n6_adj_4760), .CIN(n16113), .COUT(n16114), .S0(d6_71__N_1459[66]), 
          .S1(d6_71__N_1459[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_31 (.A0(d_tmp[64]), .B0(cout_adj_5217), .C0(n99_adj_4968), 
          .D0(n9_adj_4757), .A1(d_tmp[65]), .B1(cout_adj_5217), .C1(n96_adj_4967), 
          .D1(n8_adj_4758), .CIN(n16112), .COUT(n16113), .S0(d6_71__N_1459[64]), 
          .S1(d6_71__N_1459[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_29 (.A0(d_tmp[62]), .B0(cout_adj_5217), .C0(n105_adj_4970), 
          .D0(n11_adj_4755), .A1(d_tmp[63]), .B1(cout_adj_5217), .C1(n102_adj_4969), 
          .D1(n10_adj_4756), .CIN(n16111), .COUT(n16112), .S0(d6_71__N_1459[62]), 
          .S1(d6_71__N_1459[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_27 (.A0(d_tmp[60]), .B0(cout_adj_5217), .C0(n111_adj_4972), 
          .D0(n13_adj_4753), .A1(d_tmp[61]), .B1(cout_adj_5217), .C1(n108_adj_4971), 
          .D1(n12_adj_4754), .CIN(n16110), .COUT(n16111), .S0(d6_71__N_1459[60]), 
          .S1(d6_71__N_1459[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_25 (.A0(d_tmp[58]), .B0(cout_adj_5217), .C0(n117_adj_4974), 
          .D0(n15_adj_4751), .A1(d_tmp[59]), .B1(cout_adj_5217), .C1(n114_adj_4973), 
          .D1(n14_adj_4752), .CIN(n16109), .COUT(n16110), .S0(d6_71__N_1459[58]), 
          .S1(d6_71__N_1459[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_23 (.A0(d_tmp[56]), .B0(cout_adj_5217), .C0(n123_adj_4976), 
          .D0(n17_adj_4791), .A1(d_tmp[57]), .B1(cout_adj_5217), .C1(n120_adj_4975), 
          .D1(n16_adj_4731), .CIN(n16108), .COUT(n16109), .S0(d6_71__N_1459[56]), 
          .S1(d6_71__N_1459[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_21 (.A0(d_tmp[54]), .B0(cout_adj_5217), .C0(n129_adj_4978), 
          .D0(n19_adj_4809), .A1(d_tmp[55]), .B1(cout_adj_5217), .C1(n126_adj_4977), 
          .D1(n18_adj_4792), .CIN(n16107), .COUT(n16108), .S0(d6_71__N_1459[54]), 
          .S1(d6_71__N_1459[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_19 (.A0(d_tmp[52]), .B0(cout_adj_5217), .C0(n135_adj_4980), 
          .D0(n21_adj_4807), .A1(d_tmp[53]), .B1(cout_adj_5217), .C1(n132_adj_4979), 
          .D1(n20_adj_4808), .CIN(n16106), .COUT(n16107), .S0(d6_71__N_1459[52]), 
          .S1(d6_71__N_1459[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_17 (.A0(d_tmp[50]), .B0(cout_adj_5217), .C0(n141_adj_4982), 
          .D0(n23_adj_4805), .A1(d_tmp[51]), .B1(cout_adj_5217), .C1(n138_adj_4981), 
          .D1(n22_adj_4806), .CIN(n16105), .COUT(n16106), .S0(d6_71__N_1459[50]), 
          .S1(d6_71__N_1459[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_15 (.A0(d_tmp[48]), .B0(cout_adj_5217), .C0(n147_adj_4984), 
          .D0(n25_adj_4803), .A1(d_tmp[49]), .B1(cout_adj_5217), .C1(n144_adj_4983), 
          .D1(n24_adj_4804), .CIN(n16104), .COUT(n16105), .S0(d6_71__N_1459[48]), 
          .S1(d6_71__N_1459[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_13 (.A0(d_tmp[46]), .B0(cout_adj_5217), .C0(n153_adj_4986), 
          .D0(n27_adj_4801), .A1(d_tmp[47]), .B1(cout_adj_5217), .C1(n150_adj_4985), 
          .D1(n26_adj_4802), .CIN(n16103), .COUT(n16104), .S0(d6_71__N_1459[46]), 
          .S1(d6_71__N_1459[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_11 (.A0(d_tmp[44]), .B0(cout_adj_5217), .C0(n159_adj_4988), 
          .D0(n29_adj_4799), .A1(d_tmp[45]), .B1(cout_adj_5217), .C1(n156_adj_4987), 
          .D1(n28_adj_4800), .CIN(n16102), .COUT(n16103), .S0(d6_71__N_1459[44]), 
          .S1(d6_71__N_1459[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_9 (.A0(d_tmp[42]), .B0(cout_adj_5217), .C0(n165_adj_4990), 
          .D0(n31_adj_4797), .A1(d_tmp[43]), .B1(cout_adj_5217), .C1(n162_adj_4989), 
          .D1(n30_adj_4798), .CIN(n16101), .COUT(n16102), .S0(d6_71__N_1459[42]), 
          .S1(d6_71__N_1459[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_7 (.A0(d_tmp[40]), .B0(cout_adj_5217), .C0(n171_adj_4992), 
          .D0(n33_adj_4795), .A1(d_tmp[41]), .B1(cout_adj_5217), .C1(n168_adj_4991), 
          .D1(n32_adj_4796), .CIN(n16100), .COUT(n16101), .S0(d6_71__N_1459[40]), 
          .S1(d6_71__N_1459[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_5 (.A0(d_tmp[38]), .B0(cout_adj_5217), .C0(n177_adj_4994), 
          .D0(n35_adj_4793), .A1(d_tmp[39]), .B1(cout_adj_5217), .C1(n174_adj_4993), 
          .D1(n34_adj_4794), .CIN(n16099), .COUT(n16100), .S0(d6_71__N_1459[38]), 
          .S1(d6_71__N_1459[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_3 (.A0(d_tmp[36]), .B0(cout_adj_5217), .C0(n183_adj_4996), 
          .D0(n37_adj_4811), .A1(d_tmp[37]), .B1(cout_adj_5217), .C1(n180_adj_4995), 
          .D1(n36_adj_4810), .CIN(n16098), .COUT(n16099), .S0(d6_71__N_1459[36]), 
          .S1(d6_71__N_1459[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5217), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16098));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1460_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1460_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1460_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16094), .S0(cout_adj_5134));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1433_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1433_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_36 (.A0(d2_adj_5668[34]), .B0(d1_adj_5667[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[35]), .B1(d1_adj_5667[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16093), .COUT(n16094), .S0(d2_71__N_490_adj_5684[34]), 
          .S1(d2_71__N_490_adj_5684[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_34 (.A0(d2_adj_5668[32]), .B0(d1_adj_5667[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[33]), .B1(d1_adj_5667[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16092), .COUT(n16093), .S0(d2_71__N_490_adj_5684[32]), 
          .S1(d2_71__N_490_adj_5684[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_32 (.A0(d2_adj_5668[30]), .B0(d1_adj_5667[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[31]), .B1(d1_adj_5667[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16091), .COUT(n16092), .S0(d2_71__N_490_adj_5684[30]), 
          .S1(d2_71__N_490_adj_5684[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_30 (.A0(d2_adj_5668[28]), .B0(d1_adj_5667[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[29]), .B1(d1_adj_5667[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16090), .COUT(n16091), .S0(d2_71__N_490_adj_5684[28]), 
          .S1(d2_71__N_490_adj_5684[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_28 (.A0(d2_adj_5668[26]), .B0(d1_adj_5667[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[27]), .B1(d1_adj_5667[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16089), .COUT(n16090), .S0(d2_71__N_490_adj_5684[26]), 
          .S1(d2_71__N_490_adj_5684[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_26 (.A0(d2_adj_5668[24]), .B0(d1_adj_5667[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[25]), .B1(d1_adj_5667[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16088), .COUT(n16089), .S0(d2_71__N_490_adj_5684[24]), 
          .S1(d2_71__N_490_adj_5684[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_24 (.A0(d2_adj_5668[22]), .B0(d1_adj_5667[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[23]), .B1(d1_adj_5667[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16087), .COUT(n16088), .S0(d2_71__N_490_adj_5684[22]), 
          .S1(d2_71__N_490_adj_5684[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_22 (.A0(d2_adj_5668[20]), .B0(d1_adj_5667[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[21]), .B1(d1_adj_5667[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16086), .COUT(n16087), .S0(d2_71__N_490_adj_5684[20]), 
          .S1(d2_71__N_490_adj_5684[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_20 (.A0(d2_adj_5668[18]), .B0(d1_adj_5667[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[19]), .B1(d1_adj_5667[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16085), .COUT(n16086), .S0(d2_71__N_490_adj_5684[18]), 
          .S1(d2_71__N_490_adj_5684[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_18 (.A0(d2_adj_5668[16]), .B0(d1_adj_5667[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[17]), .B1(d1_adj_5667[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16084), .COUT(n16085), .S0(d2_71__N_490_adj_5684[16]), 
          .S1(d2_71__N_490_adj_5684[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_16 (.A0(d2_adj_5668[14]), .B0(d1_adj_5667[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[15]), .B1(d1_adj_5667[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16083), .COUT(n16084), .S0(d2_71__N_490_adj_5684[14]), 
          .S1(d2_71__N_490_adj_5684[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_14 (.A0(d2_adj_5668[12]), .B0(d1_adj_5667[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[13]), .B1(d1_adj_5667[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16082), .COUT(n16083), .S0(d2_71__N_490_adj_5684[12]), 
          .S1(d2_71__N_490_adj_5684[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_36 (.A0(d5[69]), .B0(d4[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[70]), .B1(d4[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15609), .COUT(n15610), .S0(n84_adj_5386), .S1(n81_adj_5385));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_34 (.A0(d5[67]), .B0(d4[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[68]), .B1(d4[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15608), .COUT(n15609), .S0(n90_adj_5388), .S1(n87_adj_5387));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_32 (.A0(d5[65]), .B0(d4[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[66]), .B1(d4[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15607), .COUT(n15608), .S0(n96_adj_5390), .S1(n93_adj_5389));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_30 (.A0(d5[63]), .B0(d4[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[64]), .B1(d4[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15606), .COUT(n15607), .S0(n102_adj_5392), .S1(n99_adj_5391));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_28 (.A0(d5[61]), .B0(d4[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[62]), .B1(d4[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15605), .COUT(n15606), .S0(n108_adj_5394), .S1(n105_adj_5393));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_26 (.A0(d5[59]), .B0(d4[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[60]), .B1(d4[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15604), .COUT(n15605), .S0(n114_adj_5396), .S1(n111_adj_5395));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_24 (.A0(d5[57]), .B0(d4[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[58]), .B1(d4[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15603), .COUT(n15604), .S0(n120_adj_5398), .S1(n117_adj_5397));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_22 (.A0(d5[55]), .B0(d4[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[56]), .B1(d4[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15602), .COUT(n15603), .S0(n126_adj_5400), .S1(n123_adj_5399));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_20 (.A0(d5[53]), .B0(d4[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[54]), .B1(d4[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15601), .COUT(n15602), .S0(n132_adj_5402), .S1(n129_adj_5401));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_18 (.A0(d5[51]), .B0(d4[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[52]), .B1(d4[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15600), .COUT(n15601), .S0(n138_adj_5404), .S1(n135_adj_5403));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_16 (.A0(d5[49]), .B0(d4[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[50]), .B1(d4[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15599), .COUT(n15600), .S0(n144_adj_5406), .S1(n141_adj_5405));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_14 (.A0(d5[47]), .B0(d4[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[48]), .B1(d4[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15598), .COUT(n15599), .S0(n150_adj_5408), .S1(n147_adj_5407));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_12 (.A0(d5[45]), .B0(d4[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[46]), .B1(d4[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15597), .COUT(n15598), .S0(n156_adj_5410), .S1(n153_adj_5409));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_10 (.A0(d5[43]), .B0(d4[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[44]), .B1(d4[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15596), .COUT(n15597), .S0(n162_adj_5412), .S1(n159_adj_5411));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_8 (.A0(d5[41]), .B0(d4[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[42]), .B1(d4[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15595), .COUT(n15596), .S0(n168_adj_5414), .S1(n165_adj_5413));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_6 (.A0(d5[39]), .B0(d4[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[40]), .B1(d4[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15594), .COUT(n15595), .S0(n174_adj_5416), .S1(n171_adj_5415));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_4 (.A0(d5[37]), .B0(d4[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[38]), .B1(d4[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15593), .COUT(n15594), .S0(n180_adj_5418), .S1(n177_adj_5417));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1562_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[36]), .B1(d4[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15593), .S1(n183_adj_5419));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1562_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1562_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1562_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_2.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n317), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n314), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i4 (.D(n311), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n308), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i6 (.D(n305), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n302), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i8 (.D(n299), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i9 (.D(n296), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i10 (.D(n293), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n290), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i12 (.D(n287), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i13 (.D(n284), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i14 (.D(n281), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n278), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i16 (.D(n275), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i17 (.D(n272), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i18 (.D(n269), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n266), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i20 (.D(n263), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n260), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i22 (.D(n257), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i23 (.D(n254), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n251), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i25 (.D(n248), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n245), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i27 (.D(n242), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i28 (.D(n239), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i29 (.D(n236), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n233), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i31 (.D(n230), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n227), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i33 (.D(n224), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n221), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i35 (.D(n218), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i36 (.D(n215), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i37 (.D(n212), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i38 (.D(n209_adj_4997), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i39 (.D(n206), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i40 (.D(n203), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n200), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n197), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n194), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n191), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i45 (.D(n188), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i46 (.D(n185), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n182), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i48 (.D(n179), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i49 (.D(n176), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i50 (.D(n173), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i51 (.D(n170), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n167), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i53 (.D(n164), .SP(clk_80mhz_enable_1460), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i54 (.D(n161), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i55 (.D(n158), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i56 (.D(n155), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n152), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i58 (.D(n149), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n146), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n143), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n140), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n137), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n134), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    LUT4 o_Rx_Byte_0__bdd_3_lut (.A(MYLED_0_6), .B(n17750), .C(o_Rx_Byte[3]), 
         .Z(n17521)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam o_Rx_Byte_0__bdd_3_lut.init = 16'hf6f6;
    LUT4 i3417_2_lut_2_lut (.A(o_Rx_Byte[3]), .B(n145_adj_5603), .Z(n2514)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i3417_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2445_4_lut (.A(n133), .B(n127), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12146)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2445_4_lut.init = 16'hcac0;
    LUT4 i5175_2_lut (.A(phase_inc_carrGen1[0]), .B(phase_accum_adj_5658[0]), 
         .Z(n321)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5175_2_lut.init = 16'h6666;
    LUT4 i3261_2_lut (.A(o_Rx_Byte[4]), .B(n2823), .Z(n3659)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3261_2_lut.init = 16'h4444;
    CCU2C add_3638_9 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n78_adj_5516), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n75_adj_5515), .D1(VCC_net), 
          .CIN(n16261), .COUT(n16262), .S0(n922), .S1(n921));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_9.INIT0 = 16'h9696;
    defparam add_3638_9.INIT1 = 16'h9696;
    defparam add_3638_9.INJECT1_0 = "NO";
    defparam add_3638_9.INJECT1_1 = "NO";
    LUT4 i2447_4_lut (.A(n130), .B(n124), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12148)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2447_4_lut.init = 16'hcac0;
    LUT4 i5178_2_lut (.A(MultResult2[0]), .B(MultResult1[0]), .Z(n126_adj_5178)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5178_2_lut.init = 16'h6666;
    CCU2C add_3638_7 (.A0(d_out_d_11__N_1886[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n84_adj_5518), .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n81_adj_5517), .D1(VCC_net), 
          .CIN(n16260), .COUT(n16261), .S0(n924), .S1(n923));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_7.INIT0 = 16'h9696;
    defparam add_3638_7.INIT1 = 16'h9696;
    defparam add_3638_7.INJECT1_0 = "NO";
    defparam add_3638_7.INJECT1_1 = "NO";
    LUT4 mux_325_i61_4_lut (.A(n12023), .B(n139), .C(n17625), .D(n2571), 
         .Z(n2310)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i61_4_lut.init = 16'hc0ca;
    LUT4 i2248_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n283_adj_5649), .Z(n11937)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2248_3_lut_4_lut.init = 16'hf404;
    CCU2C add_3638_5 (.A0(n90_adj_5520), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(d_out_d_11__N_1890[17]), .C1(n87_adj_5519), 
          .D1(VCC_net), .CIN(n16259), .COUT(n16260), .S0(n926), .S1(n925));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_5.INIT0 = 16'haaa0;
    defparam add_3638_5.INIT1 = 16'h9696;
    defparam add_3638_5.INJECT1_0 = "NO";
    defparam add_3638_5.INJECT1_1 = "NO";
    CCU2C add_3638_3 (.A0(d_out_d_11__N_1890[17]), .B0(ISquare[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16258), .COUT(n16259), .S1(n927));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_3.INIT0 = 16'h666a;
    defparam add_3638_3.INIT1 = 16'h555f;
    defparam add_3638_3.INJECT1_0 = "NO";
    defparam add_3638_3.INJECT1_1 = "NO";
    LUT4 i2443_4_lut (.A(n136), .B(n130_adj_5598), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12144)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2443_4_lut.init = 16'hcac0;
    LUT4 mux_325_i59_4_lut (.A(n12019), .B(n145), .C(n17625), .D(n2571), 
         .Z(n2312)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i59_4_lut.init = 16'hc0ca;
    LUT4 mux_325_i60_4_lut (.A(n12021), .B(n142), .C(n17625), .D(n2571), 
         .Z(n2311)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i60_4_lut.init = 16'hc0ca;
    CCU2C add_3638_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1890[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3638_1.INIT0 = 16'h0000;
    defparam add_3638_1.INIT1 = 16'haaaf;
    defparam add_3638_1.INJECT1_0 = "NO";
    defparam add_3638_1.INJECT1_1 = "NO";
    LUT4 i2256_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n265_adj_5643), .Z(n11945)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2256_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_325_i57_4_lut (.A(n2514), .B(n151), .C(n17625), .D(n2571), 
         .Z(n2314)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i57_4_lut.init = 16'hc0ca;
    LUT4 mux_325_i58_4_lut (.A(n2513), .B(n148), .C(n17625), .D(n2571), 
         .Z(n2313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i58_4_lut.init = 16'hcfca;
    LUT4 i3419_2_lut (.A(n142_adj_5602), .B(n17751), .Z(n2513)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3419_2_lut.init = 16'h8888;
    LUT4 mux_325_i55_4_lut (.A(n12013), .B(n157), .C(n17625), .D(n2571), 
         .Z(n2316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i55_4_lut.init = 16'hcfca;
    LUT4 mux_325_i56_4_lut (.A(n2381), .B(n154), .C(n17625), .D(n12108), 
         .Z(n2315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i56_4_lut.init = 16'hcfca;
    LUT4 i3349_2_lut (.A(n148_adj_5604), .B(n17751), .Z(n2381)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3349_2_lut.init = 16'h8888;
    CCU2C add_3634_19 (.A0(d_out_d_11__N_1886[17]), .B0(n48_adj_5422), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n45_adj_5421), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16252), .S0(n45_adj_5536), 
          .S1(d_out_d_11__N_1888[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_19.INIT0 = 16'h9995;
    defparam add_3634_19.INIT1 = 16'h9995;
    defparam add_3634_19.INJECT1_0 = "NO";
    defparam add_3634_19.INJECT1_1 = "NO";
    CCU2C add_3634_17 (.A0(d_out_d_11__N_1886[17]), .B0(n54_adj_5424), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n51_adj_5423), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16251), .COUT(n16252), .S0(n51_adj_5538), 
          .S1(n48_adj_5537));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_17.INIT0 = 16'h9995;
    defparam add_3634_17.INIT1 = 16'h9995;
    defparam add_3634_17.INJECT1_0 = "NO";
    defparam add_3634_17.INJECT1_1 = "NO";
    LUT4 i2441_4_lut (.A(n163), .B(n157_adj_5607), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12142)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2441_4_lut.init = 16'hcac0;
    LUT4 i3251_2_lut_rep_152 (.A(o_Rx_Byte[4]), .B(n2823), .Z(n17621)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3251_2_lut_rep_152.init = 16'h8888;
    LUT4 n17522_bdd_4_lut (.A(n17522), .B(n17521), .C(o_Rx_Byte[0]), .D(n17628), 
         .Z(n17618)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n17522_bdd_4_lut.init = 16'hffca;
    LUT4 mux_325_i15_4_lut (.A(n11943), .B(n277), .C(n17625), .D(n2571), 
         .Z(n2356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i15_4_lut.init = 16'hcfca;
    LUT4 i1_4_lut_4_lut_4_lut_4_lut (.A(MYLED_0_6), .B(o_Rx_Byte[0]), .C(o_Rx_Byte[4]), 
         .D(o_Rx_Byte[3]), .Z(n17027)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam i1_4_lut_4_lut_4_lut_4_lut.init = 16'h0010;
    LUT4 equal_301_i10_2_lut_2_lut (.A(MYLED_0_6), .B(o_Rx_Byte[0]), .Z(n10_adj_4732)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam equal_301_i10_2_lut_2_lut.init = 16'hdddd;
    LUT4 i6171_4_lut (.A(o_Rx_Byte[2]), .B(n16812), .C(o_Rx_Byte[3]), 
         .D(o_Rx_Byte[6]), .Z(clk_80mhz_enable_1408)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i6171_4_lut.init = 16'h0001;
    LUT4 mux_325_i16_4_lut (.A(n2555), .B(n274), .C(n17625), .D(n2571), 
         .Z(n2355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i16_4_lut.init = 16'hcfca;
    LUT4 mux_325_i54_4_lut (.A(n12011), .B(n160), .C(n17625), .D(n2571), 
         .Z(n2317)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i54_4_lut.init = 16'hc0ca;
    LUT4 i5154_2_lut (.A(d1[0]), .B(MixerOutSin[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5154_2_lut.init = 16'h6666;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i5194_2_lut (.A(d2_adj_5668[0]), .B(d1_adj_5667[0]), .Z(d2_71__N_490_adj_5684[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5194_2_lut.init = 16'h6666;
    LUT4 mux_325_i51_4_lut (.A(n2520), .B(n169), .C(n17625), .D(n2571), 
         .Z(n2320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i51_4_lut.init = 16'hcfca;
    LUT4 mux_325_i13_4_lut (.A(n2558), .B(n283), .C(n17625), .D(n2571), 
         .Z(n2358)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i13_4_lut.init = 16'hc0ca;
    LUT4 i2308_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n178_adj_5614), .Z(n11997)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2308_3_lut_4_lut.init = 16'hf404;
    LUT4 i5193_2_lut (.A(d3_adj_5669[0]), .B(d2_adj_5668[0]), .Z(d3_71__N_562_adj_5685[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5193_2_lut.init = 16'h6666;
    LUT4 i3415_2_lut (.A(n163_adj_5609), .B(o_Rx_Byte[3]), .Z(n2520)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3415_2_lut.init = 16'h8888;
    LUT4 i2433_4_lut (.A(n280), .B(n274_adj_5646), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12134)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2433_4_lut.init = 16'hcac0;
    LUT4 mux_325_i11_4_lut (.A(n11937), .B(n289), .C(n17625), .D(n2571), 
         .Z(n2360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i11_4_lut.init = 16'hcfca;
    LUT4 i5156_2_lut (.A(d1_adj_5667[0]), .B(MixerOutCos[0]), .Z(d1_71__N_418_adj_5683[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5156_2_lut.init = 16'h6666;
    LUT4 mux_325_i12_4_lut (.A(n2559), .B(n286), .C(n17625), .D(n2571), 
         .Z(n2359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i12_4_lut.init = 16'hcfca;
    LUT4 i3404_2_lut (.A(n280_adj_5648), .B(n17751), .Z(n2559)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3404_2_lut.init = 16'h8888;
    LUT4 mux_325_i9_4_lut (.A(n11933), .B(n295), .C(n17625), .D(n2571), 
         .Z(n2362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i9_4_lut.init = 16'hcfca;
    LUT4 mux_750_i22_3_lut (.A(o_Rx_Byte[2]), .B(o_Rx_Byte[4]), .C(n2823), 
         .Z(n3656)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_750_i22_3_lut.init = 16'h3a3a;
    LUT4 i2334_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n133_adj_5599), 
         .Z(n12023)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2334_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i2330_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n139_adj_5601), .Z(n12019)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2330_3_lut_4_lut.init = 16'hfb0b;
    CCU2C add_3634_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1886[17]), .C0(n60_adj_5426), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n57_adj_5425), .D1(VCC_net), .CIN(n16250), .COUT(n16251), 
          .S0(n57_adj_5540), .S1(n54_adj_5539));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_15.INIT0 = 16'h6969;
    defparam add_3634_15.INIT1 = 16'h6969;
    defparam add_3634_15.INJECT1_0 = "NO";
    defparam add_3634_15.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_37 (.A0(d4_adj_5670[70]), .B0(cout_adj_5137), 
          .C0(n81_adj_2772), .D0(d5_adj_5671[70]), .A1(d4_adj_5670[71]), 
          .B1(cout_adj_5137), .C1(n78_adj_2773), .D1(d5_adj_5671[71]), 
          .CIN(n15792), .S0(d5_71__N_706_adj_5687[70]), .S1(d5_71__N_706_adj_5687[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_37.INJECT1_1 = "NO";
    LUT4 i5190_2_lut (.A(d4_adj_5670[0]), .B(d3_adj_5669[0]), .Z(d4_71__N_634_adj_5686[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5190_2_lut.init = 16'h6666;
    LUT4 i5187_2_lut (.A(d5_adj_5671[0]), .B(d4_adj_5670[0]), .Z(d5_71__N_706_adj_5687[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5187_2_lut.init = 16'h6666;
    CCU2C add_3634_13 (.A0(d_out_d_11__N_1886[17]), .B0(n66_adj_5428), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n63_adj_5427), .D1(VCC_net), .CIN(n16249), .COUT(n16250), 
          .S0(n63_adj_5542), .S1(n60_adj_5541));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_13.INIT0 = 16'h9995;
    defparam add_3634_13.INIT1 = 16'h6969;
    defparam add_3634_13.INJECT1_0 = "NO";
    defparam add_3634_13.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_35 (.A0(d4_adj_5670[68]), .B0(cout_adj_5137), 
          .C0(n87_adj_2770), .D0(d5_adj_5671[68]), .A1(d4_adj_5670[69]), 
          .B1(cout_adj_5137), .C1(n84_adj_2771), .D1(d5_adj_5671[69]), 
          .CIN(n15791), .COUT(n15792), .S0(d5_71__N_706_adj_5687[68]), 
          .S1(d5_71__N_706_adj_5687[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_33 (.A0(d4_adj_5670[66]), .B0(cout_adj_5137), 
          .C0(n93), .D0(d5_adj_5671[66]), .A1(d4_adj_5670[67]), .B1(cout_adj_5137), 
          .C1(n90_adj_2769), .D1(d5_adj_5671[67]), .CIN(n15790), .COUT(n15791), 
          .S0(d5_71__N_706_adj_5687[66]), .S1(d5_71__N_706_adj_5687[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_12 (.A0(d2_adj_5668[10]), .B0(d1_adj_5667[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[11]), .B1(d1_adj_5667[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16081), .COUT(n16082), .S0(d2_71__N_490_adj_5684[10]), 
          .S1(d2_71__N_490_adj_5684[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_12.INJECT1_1 = "NO";
    CCU2C add_3634_11 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n72_adj_5430), .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), 
          .B1(n17635), .C1(n69_adj_5429), .D1(VCC_net), .CIN(n16248), 
          .COUT(n16249), .S0(n69_adj_5544), .S1(n66_adj_5543));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_11.INIT0 = 16'h9696;
    defparam add_3634_11.INIT1 = 16'h6969;
    defparam add_3634_11.INJECT1_0 = "NO";
    defparam add_3634_11.INJECT1_1 = "NO";
    CCU2C add_3634_9 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n78_adj_5432), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n75_adj_5431), .D1(VCC_net), 
          .CIN(n16247), .COUT(n16248), .S0(n75_adj_5546), .S1(n72_adj_5545));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_9.INIT0 = 16'h9696;
    defparam add_3634_9.INIT1 = 16'h9696;
    defparam add_3634_9.INJECT1_0 = "NO";
    defparam add_3634_9.INJECT1_1 = "NO";
    CCU2C add_3634_7 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n84_adj_5434), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n81_adj_5433), .D1(VCC_net), 
          .CIN(n16246), .COUT(n16247), .S0(n81_adj_5548), .S1(n78_adj_5547));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_7.INIT0 = 16'h9696;
    defparam add_3634_7.INIT1 = 16'h9696;
    defparam add_3634_7.INJECT1_0 = "NO";
    defparam add_3634_7.INJECT1_1 = "NO";
    CCU2C add_3634_5 (.A0(n90_adj_5436), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(d_out_d_11__N_1886[17]), .C1(n87_adj_5435), 
          .D1(VCC_net), .CIN(n16245), .COUT(n16246), .S0(n87_adj_5550), 
          .S1(n84_adj_5549));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_5.INIT0 = 16'haaa0;
    defparam add_3634_5.INIT1 = 16'h9696;
    defparam add_3634_5.INJECT1_0 = "NO";
    defparam add_3634_5.INJECT1_1 = "NO";
    CCU2C add_3634_3 (.A0(d_out_d_11__N_1886[17]), .B0(ISquare[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16244), .COUT(n16245), .S1(n90_adj_5551));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_3.INIT0 = 16'h666a;
    defparam add_3634_3.INIT1 = 16'h555f;
    defparam add_3634_3.INJECT1_0 = "NO";
    defparam add_3634_3.INJECT1_1 = "NO";
    CCU2C add_3634_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16244));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3634_1.INIT0 = 16'h0000;
    defparam add_3634_1.INIT1 = 16'haaaf;
    defparam add_3634_1.INJECT1_0 = "NO";
    defparam add_3634_1.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_10 (.A0(d2_adj_5668[8]), .B0(d1_adj_5667[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[9]), .B1(d1_adj_5667[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16080), .COUT(n16081), .S0(d2_71__N_490_adj_5684[8]), 
          .S1(d2_71__N_490_adj_5684[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_10.INJECT1_1 = "NO";
    CCU2C add_3636_19 (.A0(d_out_d_11__N_1879), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1879), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16238), .S0(n45_adj_5489), 
          .S1(d_out_d_11__N_1882[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_19.INIT0 = 16'h666a;
    defparam add_3636_19.INIT1 = 16'h666a;
    defparam add_3636_19.INJECT1_0 = "NO";
    defparam add_3636_19.INJECT1_1 = "NO";
    CCU2C add_3636_17 (.A0(d_out_d_11__N_1880[17]), .B0(n54_adj_5256), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n51_adj_5255), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16237), .COUT(n16238), .S0(n51_adj_5491), 
          .S1(n48_adj_5490));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_17.INIT0 = 16'h9995;
    defparam add_3636_17.INIT1 = 16'h9995;
    defparam add_3636_17.INJECT1_0 = "NO";
    defparam add_3636_17.INJECT1_1 = "NO";
    CCU2C add_3636_15 (.A0(d_out_d_11__N_1880[17]), .B0(n60_adj_5258), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n57_adj_5257), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16236), .COUT(n16237), .S0(n57_adj_5493), 
          .S1(n54_adj_5492));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_15.INIT0 = 16'h9995;
    defparam add_3636_15.INIT1 = 16'h9995;
    defparam add_3636_15.INJECT1_0 = "NO";
    defparam add_3636_15.INJECT1_1 = "NO";
    CCU2C add_3636_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n66_adj_5260), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n63_adj_5259), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16235), .COUT(n16236), .S0(n63_adj_5495), 
          .S1(n60_adj_5494));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_13.INIT0 = 16'h6969;
    defparam add_3636_13.INIT1 = 16'h9995;
    defparam add_3636_13.INJECT1_0 = "NO";
    defparam add_3636_13.INJECT1_1 = "NO";
    CCU2C add_3636_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n72_adj_5262), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1880[17]), 
          .C1(n69_adj_5261), .D1(VCC_net), .CIN(n16234), .COUT(n16235), 
          .S0(n69_adj_5497), .S1(n66_adj_5496));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_11.INIT0 = 16'h6969;
    defparam add_3636_11.INIT1 = 16'h6969;
    defparam add_3636_11.INJECT1_0 = "NO";
    defparam add_3636_11.INJECT1_1 = "NO";
    CCU2C add_3636_9 (.A0(d_out_d_11__N_1880[17]), .B0(n17635), .C0(n78_adj_5264), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n75_adj_5263), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16233), .COUT(n16234), .S0(n75_adj_5499), 
          .S1(n72_adj_5498));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_9.INIT0 = 16'h6969;
    defparam add_3636_9.INIT1 = 16'h9995;
    defparam add_3636_9.INJECT1_0 = "NO";
    defparam add_3636_9.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_11 (.A0(d6[44]), .B0(cout_adj_5341), .C0(n159_adj_4952), 
          .D0(n29_adj_4706), .A1(d6[45]), .B1(cout_adj_5341), .C1(n156_adj_4951), 
          .D1(n28_adj_4707), .CIN(n16006), .COUT(n16007), .S0(d7_71__N_1531[44]), 
          .S1(d7_71__N_1531[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_11.INJECT1_1 = "NO";
    CCU2C add_3636_7 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(n84_adj_5266), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1880[17]), .C1(n81_adj_5265), .D1(VCC_net), 
          .CIN(n16232), .COUT(n16233), .S0(n81_adj_5501), .S1(n78_adj_5500));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_7.INIT0 = 16'h9696;
    defparam add_3636_7.INIT1 = 16'h9696;
    defparam add_3636_7.INJECT1_0 = "NO";
    defparam add_3636_7.INJECT1_1 = "NO";
    CCU2C add_3636_5 (.A0(n90_adj_5268), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1880[17]), .C1(n87_adj_5267), 
          .D1(VCC_net), .CIN(n16231), .COUT(n16232), .S0(n87_adj_5503), 
          .S1(n84_adj_5502));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_5.INIT0 = 16'haaa0;
    defparam add_3636_5.INIT1 = 16'h9696;
    defparam add_3636_5.INJECT1_0 = "NO";
    defparam add_3636_5.INJECT1_1 = "NO";
    LUT4 mux_325_i10_4_lut (.A(n11935), .B(n292), .C(n17625), .D(n2571), 
         .Z(n2361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i10_4_lut.init = 16'hcfca;
    LUT4 i2431_4_lut (.A(n301), .B(n295_adj_5653), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2431_4_lut.init = 16'hcacf;
    LUT4 mux_325_i8_4_lut (.A(n2563), .B(n298), .C(n17625), .D(n2571), 
         .Z(n2363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i8_4_lut.init = 16'hcfca;
    LUT4 mux_325_i5_4_lut (.A(n11927), .B(n307), .C(n17625), .D(n2571), 
         .Z(n2366)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i5_4_lut.init = 16'hc0ca;
    LUT4 i3402_1_lut_2_lut (.A(o_Rx_Byte[4]), .B(n2823), .Z(n3676)) /* synthesis lut_function=(!(A (B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3402_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_325_i52_4_lut (.A(n12007), .B(n166), .C(n17625), .D(n2571), 
         .Z(n2319)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i52_4_lut.init = 16'hc0ca;
    CCU2C add_3636_3 (.A0(d_out_d_11__N_1880[17]), .B0(ISquare[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16230), .COUT(n16231), .S1(n90_adj_5504));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_3.INIT0 = 16'h666a;
    defparam add_3636_3.INIT1 = 16'h555f;
    defparam add_3636_3.INJECT1_0 = "NO";
    defparam add_3636_3.INJECT1_1 = "NO";
    CCU2C add_3636_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16230));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam add_3636_1.INIT0 = 16'h0000;
    defparam add_3636_1.INIT1 = 16'haaaf;
    defparam add_3636_1.INJECT1_0 = "NO";
    defparam add_3636_1.INJECT1_1 = "NO";
    LUT4 i6154_4_lut (.A(n17784), .B(o_Rx_Byte[3]), .C(n13169), .D(n17629), 
         .Z(clk_80mhz_enable_45)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;
    defparam i6154_4_lut.init = 16'ha0a2;
    LUT4 mux_325_i6_4_lut (.A(n11929), .B(n304), .C(n17625), .D(n2571), 
         .Z(n2365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i6_4_lut.init = 16'hcfca;
    LUT4 i2298_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n199_adj_5621), .Z(n11987)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2298_3_lut_4_lut.init = 16'hf404;
    LUT4 i2268_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n244_adj_5636), 
         .Z(n11957)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2268_3_lut_4_lut.init = 16'hf404;
    LUT4 i6166_4_lut (.A(n16740), .B(n17632), .C(n17648), .D(n17449), 
         .Z(clk_80mhz_enable_1470)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i6166_4_lut.init = 16'h3032;
    LUT4 i2332_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n136_adj_5600), .Z(n12021)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2332_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i15_3_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[3]), .C(o_Rx_Byte[0]), 
         .Z(n16740)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i15_3_lut.init = 16'h3636;
    LUT4 mux_325_i49_4_lut (.A(n12003), .B(n175), .C(n17625), .D(n2571), 
         .Z(n2322)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i49_4_lut.init = 16'hc0ca;
    LUT4 i2324_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n151_adj_5605), .Z(n12013)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2324_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_325_i50_4_lut (.A(n2387), .B(n172), .C(n17625), .D(n12108), 
         .Z(n2321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i50_4_lut.init = 16'hcfca;
    LUT4 i3348_2_lut (.A(n166_adj_5610), .B(n17751), .Z(n2387)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3348_2_lut.init = 16'h8888;
    LUT4 i3266_rep_84_2_lut (.A(o_Rx_Byte[2]), .B(MYLED_0_6), .Z(n17449)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3266_rep_84_2_lut.init = 16'heeee;
    LUT4 i2284_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n220_adj_5628), .Z(n11973)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2284_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_325_i47_4_lut (.A(n11999), .B(n181), .C(n17625), .D(n2571), 
         .Z(n2324)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i47_4_lut.init = 16'hc0ca;
    LUT4 i2294_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n205_adj_5623), .Z(n11983)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2294_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_325_i3_4_lut (.A(o_Rx_Byte[3]), .B(n313), .C(n17625), .D(n17631), 
         .Z(n2368)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i3_4_lut.init = 16'hc0c5;
    LUT4 i2300_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n196_adj_5620), 
         .Z(n11989)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2300_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_325_i48_4_lut (.A(n12001), .B(n178), .C(n17625), .D(n2571), 
         .Z(n2323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i48_4_lut.init = 16'hcfca;
    LUT4 mux_325_i2_4_lut (.A(n12511), .B(n316), .C(n17625), .D(n2571), 
         .Z(n2369)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i2_4_lut.init = 16'hcfc5;
    LUT4 mux_325_i45_4_lut (.A(n2392), .B(n187), .C(n17625), .D(n12108), 
         .Z(n2326)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i45_4_lut.init = 16'hc0ca;
    LUT4 i2312_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n172_adj_5612), .Z(n12001)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2312_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i6159_4_lut (.A(n12378), .B(o_Rx_Byte[2]), .C(n17573), .D(n17633), 
         .Z(n13169)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i6159_4_lut.init = 16'h575f;
    LUT4 i2278_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n229_adj_5631), 
         .Z(n11967)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2278_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_325_i46_4_lut (.A(n11997), .B(n184), .C(n17625), .D(n2571), 
         .Z(n2325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i46_4_lut.init = 16'hcfca;
    LUT4 i2306_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n184_adj_5616), .Z(n11995)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2306_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_750_i3_3_lut_rep_153 (.A(o_Rx_Byte[2]), .B(o_Rx_Byte[4]), .C(n2823), 
         .Z(n17622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_750_i3_3_lut_rep_153.init = 16'hcaca;
    FD1S3AX o_Rx_Byte_i3_rep_175 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(n17751));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i3_rep_175.GSR = "ENABLED";
    CCU2C _add_1_1490_add_4_31 (.A0(d4_adj_5670[64]), .B0(cout_adj_5137), 
          .C0(n99), .D0(d5_adj_5671[64]), .A1(d4_adj_5670[65]), .B1(cout_adj_5137), 
          .C1(n96), .D1(d5_adj_5671[65]), .CIN(n15789), .COUT(n15790), 
          .S0(d5_71__N_706_adj_5687[64]), .S1(d5_71__N_706_adj_5687[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(70[13:20])
    defparam _add_1_1490_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1490_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1490_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_8 (.A0(d2_adj_5668[6]), .B0(d1_adj_5667[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[7]), .B1(d1_adj_5667[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16079), .COUT(n16080), .S0(d2_71__N_490_adj_5684[6]), 
          .S1(d2_71__N_490_adj_5684[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_23 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n123_adj_5105), .D0(d1[56]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n120_adj_5104), .D1(d1[57]), .CIN(n15860), .COUT(n15861), 
          .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_6 (.A0(d2_adj_5668[4]), .B0(d1_adj_5667[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[5]), .B1(d1_adj_5667[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16078), .COUT(n16079), .S0(d2_71__N_490_adj_5684[4]), 
          .S1(d2_71__N_490_adj_5684[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_4 (.A0(d2_adj_5668[2]), .B0(d1_adj_5667[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[3]), .B1(d1_adj_5667[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16077), .COUT(n16078), .S0(d2_71__N_490_adj_5684[2]), 
          .S1(d2_71__N_490_adj_5684[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_9 (.A0(d6[42]), .B0(cout_adj_5341), .C0(n165_adj_4954), 
          .D0(n31_adj_4704), .A1(d6[43]), .B1(cout_adj_5341), .C1(n162_adj_4953), 
          .D1(n30_adj_4705), .CIN(n16005), .COUT(n16006), .S0(d7_71__N_1531[42]), 
          .S1(d7_71__N_1531[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_2 (.A0(d2_adj_5668[0]), .B0(d1_adj_5667[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5668[1]), .B1(d1_adj_5667[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16077), .S1(d2_71__N_490_adj_5684[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(64[13:20])
    defparam _add_1_1433_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1433_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_6 (.A0(d_d_tmp[3]), .B0(d_tmp[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[4]), .B1(d_tmp[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16022), .COUT(n16023), .S0(d6_71__N_1459[3]), 
          .S1(d6_71__N_1459[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16075), .S0(cout_adj_5135));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1436_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1436_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_7 (.A0(d6[40]), .B0(cout_adj_5341), .C0(n171_adj_4956), 
          .D0(n33_adj_4702), .A1(d6[41]), .B1(cout_adj_5341), .C1(n168_adj_4955), 
          .D1(n32_adj_4703), .CIN(n16004), .COUT(n16005), .S0(d7_71__N_1531[40]), 
          .S1(d7_71__N_1531[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_36 (.A0(d3_adj_5669[34]), .B0(d2_adj_5668[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[35]), .B1(d2_adj_5668[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16074), .COUT(n16075), .S0(d3_71__N_562_adj_5685[34]), 
          .S1(d3_71__N_562_adj_5685[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_34 (.A0(d3_adj_5669[32]), .B0(d2_adj_5668[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[33]), .B1(d2_adj_5668[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16073), .COUT(n16074), .S0(d3_71__N_562_adj_5685[32]), 
          .S1(d3_71__N_562_adj_5685[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_32 (.A0(d3_adj_5669[30]), .B0(d2_adj_5668[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[31]), .B1(d2_adj_5668[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16072), .COUT(n16073), .S0(d3_71__N_562_adj_5685[30]), 
          .S1(d3_71__N_562_adj_5685[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_30 (.A0(d3_adj_5669[28]), .B0(d2_adj_5668[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[29]), .B1(d2_adj_5668[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16071), .COUT(n16072), .S0(d3_71__N_562_adj_5685[28]), 
          .S1(d3_71__N_562_adj_5685[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_28 (.A0(d3_adj_5669[26]), .B0(d2_adj_5668[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[27]), .B1(d2_adj_5668[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16070), .COUT(n16071), .S0(d3_71__N_562_adj_5685[26]), 
          .S1(d3_71__N_562_adj_5685[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_21 (.A0(MixerOutSin[11]), .B0(cout_adj_4999), 
          .C0(n129_adj_5107), .D0(d1[54]), .A1(MixerOutSin[11]), .B1(cout_adj_4999), 
          .C1(n126_adj_5106), .D1(d1[55]), .CIN(n15859), .COUT(n15860), 
          .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(62[13:22])
    defparam _add_1_1448_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_26 (.A0(d3_adj_5669[24]), .B0(d2_adj_5668[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[25]), .B1(d2_adj_5668[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16069), .COUT(n16070), .S0(d3_71__N_562_adj_5685[24]), 
          .S1(d3_71__N_562_adj_5685[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_24 (.A0(d3_adj_5669[22]), .B0(d2_adj_5668[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[23]), .B1(d2_adj_5668[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16068), .COUT(n16069), .S0(d3_71__N_562_adj_5685[22]), 
          .S1(d3_71__N_562_adj_5685[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_4 (.A0(d_d_tmp[1]), .B0(d_tmp[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[2]), .B1(d_tmp[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16021), .COUT(n16022), .S0(d6_71__N_1459[1]), 
          .S1(d6_71__N_1459[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_22 (.A0(d3_adj_5669[20]), .B0(d2_adj_5668[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[21]), .B1(d2_adj_5668[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16067), .COUT(n16068), .S0(d3_71__N_562_adj_5685[20]), 
          .S1(d3_71__N_562_adj_5685[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_22.INJECT1_1 = "NO";
    LUT4 i2292_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n208_adj_5624), 
         .Z(n11981)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2292_3_lut_4_lut.init = 16'hf404;
    LUT4 i2238_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n301_adj_5655), .Z(n11927)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2238_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1436_add_4_20 (.A0(d3_adj_5669[18]), .B0(d2_adj_5668[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[19]), .B1(d2_adj_5668[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16066), .COUT(n16067), .S0(d3_71__N_562_adj_5685[18]), 
          .S1(d3_71__N_562_adj_5685[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_18 (.A0(d3_adj_5669[16]), .B0(d2_adj_5668[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[17]), .B1(d2_adj_5668[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16065), .COUT(n16066), .S0(d3_71__N_562_adj_5685[16]), 
          .S1(d3_71__N_562_adj_5685[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_5 (.A0(d6[38]), .B0(cout_adj_5341), .C0(n177_adj_4958), 
          .D0(n35_adj_4700), .A1(d6[39]), .B1(cout_adj_5341), .C1(n174_adj_4957), 
          .D1(n34_adj_4701), .CIN(n16003), .COUT(n16004), .S0(d7_71__N_1531[38]), 
          .S1(d7_71__N_1531[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[0]), .B1(d_tmp[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16021), .S1(d6_71__N_1459[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1520_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_2.INJECT1_1 = "NO";
    PLL PLL1 (.osc_clk_c(osc_clk_c), .clk_80mhz(clk_80mhz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(124[5] 127[2])
    CCU2C _add_1_1463_add_4_37 (.A0(d6[70]), .B0(cout_adj_5341), .C0(n81_adj_4926), 
          .D0(n3_adj_4568), .A1(d6[71]), .B1(cout_adj_5341), .C1(n78_adj_4925), 
          .D1(n2_adj_4569), .CIN(n16019), .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_35 (.A0(d6[68]), .B0(cout_adj_5341), .C0(n87_adj_4928), 
          .D0(n5_adj_4730), .A1(d6[69]), .B1(cout_adj_5341), .C1(n84_adj_4927), 
          .D1(n4_adj_4567), .CIN(n16018), .COUT(n16019), .S0(d7_71__N_1531[68]), 
          .S1(d7_71__N_1531[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_33 (.A0(d6[66]), .B0(cout_adj_5341), .C0(n93_adj_4930), 
          .D0(n7_adj_4728), .A1(d6[67]), .B1(cout_adj_5341), .C1(n90_adj_4929), 
          .D1(n6_adj_4729), .CIN(n16017), .COUT(n16018), .S0(d7_71__N_1531[66]), 
          .S1(d7_71__N_1531[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_31 (.A0(d6[64]), .B0(cout_adj_5341), .C0(n99_adj_4932), 
          .D0(n9_adj_4726), .A1(d6[65]), .B1(cout_adj_5341), .C1(n96_adj_4931), 
          .D1(n8_adj_4727), .CIN(n16016), .COUT(n16017), .S0(d7_71__N_1531[64]), 
          .S1(d7_71__N_1531[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_31.INJECT1_1 = "NO";
    LUT4 mux_325_i43_4_lut (.A(n11993), .B(n193), .C(n17625), .D(n2571), 
         .Z(n2328)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i43_4_lut.init = 16'hc0ca;
    LUT4 i2286_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n217_adj_5627), .Z(n11975)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2286_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1463_add_4_29 (.A0(d6[62]), .B0(cout_adj_5341), .C0(n105_adj_4934), 
          .D0(n11_adj_4724), .A1(d6[63]), .B1(cout_adj_5341), .C1(n102_adj_4933), 
          .D1(n10_adj_4725), .CIN(n16015), .COUT(n16016), .S0(d7_71__N_1531[62]), 
          .S1(d7_71__N_1531[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_27 (.A0(d6[60]), .B0(cout_adj_5341), .C0(n111_adj_4936), 
          .D0(n13_adj_4722), .A1(d6[61]), .B1(cout_adj_5341), .C1(n108_adj_4935), 
          .D1(n12_adj_4723), .CIN(n16014), .COUT(n16015), .S0(d7_71__N_1531[60]), 
          .S1(d7_71__N_1531[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_25 (.A0(d6[58]), .B0(cout_adj_5341), .C0(n117_adj_4938), 
          .D0(n15_adj_4720), .A1(d6[59]), .B1(cout_adj_5341), .C1(n114_adj_4937), 
          .D1(n14_adj_4721), .CIN(n16013), .COUT(n16014), .S0(d7_71__N_1531[58]), 
          .S1(d7_71__N_1531[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_25.INJECT1_1 = "NO";
    LUT4 i2288_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n214_adj_5626), .Z(n11977)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2288_3_lut_4_lut.init = 16'hfb0b;
    CCU2C ISquare_add_4_16 (.A0(MultResult2[14]), .B0(MultResult1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[15]), .B1(MultResult1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15801), .COUT(n15802), .S0(n84_adj_5164), 
          .S1(n81_adj_5163));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_16.INIT0 = 16'h666a;
    defparam ISquare_add_4_16.INIT1 = 16'h666a;
    defparam ISquare_add_4_16.INJECT1_0 = "NO";
    defparam ISquare_add_4_16.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_18 (.A0(MultResult2[16]), .B0(MultResult1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[17]), .B1(MultResult1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15802), .COUT(n15803), .S0(n78_adj_5162), 
          .S1(n75_adj_5161));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(92[16:41])
    defparam ISquare_add_4_18.INIT0 = 16'h666a;
    defparam ISquare_add_4_18.INIT1 = 16'h666a;
    defparam ISquare_add_4_18.INJECT1_0 = "NO";
    defparam ISquare_add_4_18.INJECT1_1 = "NO";
    LUT4 i2270_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n241_adj_5635), .Z(n11959)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2270_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_4_lut (.A(o_Rx_Byte[7]), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[6]), 
         .D(o_Rx_DV), .Z(n12378)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h4000;
    LUT4 i2322_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n154_adj_5606), 
         .Z(n12011)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2322_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_325_i44_4_lut (.A(n11995), .B(n190), .C(n17625), .D(n2571), 
         .Z(n2327)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i44_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1619_add_4_4 (.A0(d_d9[1]), .B0(d9[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[2]), .B1(d9[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14899), .COUT(n14900));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam _add_1_1619_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1619_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1619_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1619_add_4_4.INJECT1_1 = "NO";
    LUT4 mux_325_i41_4_lut (.A(n2530), .B(n199), .C(n17625), .D(n2571), 
         .Z(n2330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i41_4_lut.init = 16'hcfca;
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 i2439_4_lut (.A(n196), .B(n190_adj_5618), .C(o_Rx_Byte[3]), .D(n17629), 
         .Z(n12140)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2439_4_lut.init = 16'hcac0;
    CCU2C _add_1_1436_add_4_16 (.A0(d3_adj_5669[14]), .B0(d2_adj_5668[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[15]), .B1(d2_adj_5668[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16064), .COUT(n16065), .S0(d3_71__N_562_adj_5685[14]), 
          .S1(d3_71__N_562_adj_5685[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_16.INJECT1_1 = "NO";
    LUT4 i2314_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n169_adj_5611), .Z(n12003)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2314_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_325_i39_4_lut (.A(n11987), .B(n205), .C(n17625), .D(n2571), 
         .Z(n2332)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i39_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1436_add_4_14 (.A0(d3_adj_5669[12]), .B0(d2_adj_5668[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[13]), .B1(d2_adj_5668[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16063), .COUT(n16064), .S0(d3_71__N_562_adj_5685[12]), 
          .S1(d3_71__N_562_adj_5685[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_14.INJECT1_1 = "NO";
    LUT4 mux_325_i40_4_lut (.A(n11989), .B(n202), .C(n17625), .D(n2571), 
         .Z(n2331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i40_4_lut.init = 16'hcfca;
    CCU2C _add_1_1436_add_4_12 (.A0(d3_adj_5669[10]), .B0(d2_adj_5668[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[11]), .B1(d2_adj_5668[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16062), .COUT(n16063), .S0(d3_71__N_562_adj_5685[10]), 
          .S1(d3_71__N_562_adj_5685[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_12.INJECT1_1 = "NO";
    LUT4 mux_325_i37_4_lut (.A(n11983), .B(n211), .C(n17625), .D(n2571), 
         .Z(n2334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i37_4_lut.init = 16'hcfca;
    CCU2C _add_1_1436_add_4_10 (.A0(d3_adj_5669[8]), .B0(d2_adj_5668[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[9]), .B1(d2_adj_5668[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16061), .COUT(n16062), .S0(d3_71__N_562_adj_5685[8]), 
          .S1(d3_71__N_562_adj_5685[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_10.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i1 (.D(n320), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    LUT4 i2310_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n175_adj_5613), .Z(n11999)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2310_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_325_i38_4_lut (.A(n11985), .B(n208), .C(n17625), .D(n2571), 
         .Z(n2333)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i38_4_lut.init = 16'hc0ca;
    LUT4 i3252_2_lut (.A(o_Rx_Byte[4]), .B(n2823), .Z(n3677)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i3252_2_lut.init = 16'hbbbb;
    LUT4 mux_325_i35_4_lut (.A(n11979), .B(n217), .C(n17625), .D(n2571), 
         .Z(n2336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i35_4_lut.init = 16'hcfca;
    LUT4 mux_325_i36_4_lut (.A(n11981), .B(n214), .C(n17625), .D(n2571), 
         .Z(n2335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i36_4_lut.init = 16'hcfca;
    LUT4 i2304_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n187_adj_5617), 
         .Z(n11993)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2304_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_325_i33_4_lut (.A(n11975), .B(n223), .C(n17625), .D(n2571), 
         .Z(n2338)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i33_4_lut.init = 16'hc0ca;
    LUT4 i2006_1_lut_3_lut (.A(o_Rx_Byte[2]), .B(o_Rx_Byte[4]), .C(n2823), 
         .Z(n11690)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2006_1_lut_3_lut.init = 16'h3535;
    LUT4 mux_325_i34_4_lut (.A(n11977), .B(n220), .C(n17625), .D(n2571), 
         .Z(n2337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i34_4_lut.init = 16'hcfca;
    LUT4 i2296_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n202_adj_5622), .Z(n11985)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2296_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_325_i31_4_lut (.A(n11971), .B(n229), .C(n17625), .D(n2571), 
         .Z(n2340)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i31_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1436_add_4_8 (.A0(d3_adj_5669[6]), .B0(d2_adj_5668[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[7]), .B1(d2_adj_5668[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16060), .COUT(n16061), .S0(d3_71__N_562_adj_5685[6]), 
          .S1(d3_71__N_562_adj_5685[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_8.INJECT1_1 = "NO";
    LUT4 mux_325_i32_4_lut (.A(n11973), .B(n226), .C(n17625), .D(n2571), 
         .Z(n2339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i32_4_lut.init = 16'hcfca;
    LUT4 mux_750_i2_3_lut (.A(o_Rx_Byte[2]), .B(o_Rx_Byte[4]), .C(n2823), 
         .Z(n3691)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_750_i2_3_lut.init = 16'hc5c5;
    LUT4 i2318_3_lut_4_lut (.A(n17750), .B(n17630), .C(n17751), .D(n160_adj_5608), 
         .Z(n12007)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2318_3_lut_4_lut.init = 16'hf404;
    LUT4 i2290_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n211_adj_5625), .Z(n11979)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2290_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_325_i29_4_lut (.A(n11967), .B(n235), .C(n17625), .D(n2571), 
         .Z(n2342)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i29_4_lut.init = 16'hc0ca;
    LUT4 i2282_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n223_adj_5629), .Z(n11971)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2282_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1436_add_4_6 (.A0(d3_adj_5669[4]), .B0(d2_adj_5668[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[5]), .B1(d2_adj_5668[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16059), .COUT(n16060), .S0(d3_71__N_562_adj_5685[4]), 
          .S1(d3_71__N_562_adj_5685[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_6.INJECT1_1 = "NO";
    LUT4 mux_325_i30_4_lut (.A(n2541), .B(n232), .C(n17625), .D(n2571), 
         .Z(n2341)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i30_4_lut.init = 16'hc0ca;
    LUT4 i2274_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n235_adj_5633), .Z(n11963)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2274_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_325_i27_4_lut (.A(n11963), .B(n241), .C(n17625), .D(n2571), 
         .Z(n2344)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i27_4_lut.init = 16'hc0ca;
    LUT4 i1_3_lut_rep_164_3_lut (.A(o_Rx_Byte[0]), .B(MYLED_0_6), .C(o_Rx_Byte[4]), 
         .Z(n17633)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_3_lut_rep_164_3_lut.init = 16'h0404;
    CCU2C _add_1_1436_add_4_4 (.A0(d3_adj_5669[2]), .B0(d2_adj_5668[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[3]), .B1(d2_adj_5668[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16058), .COUT(n16059), .S0(d3_71__N_562_adj_5685[2]), 
          .S1(d3_71__N_562_adj_5685[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_2 (.A0(d3_adj_5669[0]), .B0(d2_adj_5668[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5669[1]), .B1(d2_adj_5668[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16058), .S1(d3_71__N_562_adj_5685[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(66[13:20])
    defparam _add_1_1436_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1436_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_2.INJECT1_1 = "NO";
    LUT4 mux_325_i28_4_lut (.A(n11965), .B(n238), .C(n17625), .D(n2571), 
         .Z(n2343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i28_4_lut.init = 16'hcfca;
    LUT4 i2276_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n17630), .C(n17751), 
         .D(n232_adj_5632), .Z(n11965)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2276_3_lut_4_lut.init = 16'hf707;
    LUT4 i1_2_lut_rep_161_4_lut_4_lut (.A(o_Rx_Byte[0]), .B(n12378), .C(MYLED_0_6), 
         .D(o_Rx_Byte[4]), .Z(n17630)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_2_lut_rep_161_4_lut_4_lut.init = 16'h0040;
    CCU2C _add_1_1559_add_4_38 (.A0(d4[71]), .B0(d3[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16056), .S0(n78_adj_5342));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1559_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_38.INJECT1_1 = "NO";
    \CIC(width=72,decimation_ratio=4096)  CIC1Sin (.d_tmp({d_tmp}), .clk_80mhz(clk_80mhz), 
            .d5({d5}), .d_d_tmp({d_d_tmp}), .d_d7({d_d7}), .n29(n29), 
            .n28(n28), .d2({d2}), .d2_71__N_490({d2_71__N_490}), .d3({d3}), 
            .d3_71__N_562({d3_71__N_562}), .n7(n7_adj_4759), .d4({d4}), 
            .d4_71__N_634({d4_71__N_634}), .d5_71__N_706({d5_71__N_706}), 
            .d6({d6}), .d6_71__N_1459({d6_71__N_1459}), .d_d6({d_d6}), 
            .CIC1_out_clkSin(CIC1_out_clkSin), .d7({d7}), .d7_71__N_1531({d7_71__N_1531}), 
            .d8({d8}), .d8_71__N_1603({d8_71__N_1603}), .d_d8({d_d8}), 
            .d9({d9}), .d9_71__N_1675({d9_71__N_1675}), .d_d9({d_d9}), 
            .n6(n6_adj_4760), .\CIC1_outSin[0] (CIC1_outSin[0]), .d1({d1}), 
            .d1_71__N_418({d1_71__N_418}), .count({count}), .n9(n9_adj_4757), 
            .n8(n8_adj_4758), .n11(n11_adj_4755), .n10(n10_adj_4756), 
            .n13(n13_adj_4753), .n12(n12_adj_4754), .n31(n31), .n30(n30), 
            .n33(n33_adj_4697), .n15(n15_adj_4751), .n14(n14_adj_4752), 
            .n17(n17_adj_4791), .n16(n16_adj_4731), .n19(n19_adj_4809), 
            .n18(n18_adj_4792), .n32(n32), .n5(n5_adj_4832), .n4(n4_adj_4833), 
            .n35(n35_adj_4695), .n7_adj_115(n7_adj_4830), .n21(n21_adj_4807), 
            .n20(n20_adj_4808), .n23(n23_adj_4805), .n22(n22_adj_4806), 
            .n25(n25_adj_4803), .n24(n24_adj_4781), .n27(n27_adj_4778), 
            .n34(n34_adj_4696), .\CICGain[1] (CICGain[1]), .\CICGain[0] (CICGain[0]), 
            .\d10[66] (d10_adj_5680[66]), .\d10[67] (d10_adj_5680[67]), 
            .n26(n26_adj_4779), .n29_adj_116(n29_adj_4776), .\d10[69] (d10_adj_5680[69]), 
            .\d10[68] (d10_adj_5680[68]), .n28_adj_117(n28_adj_4777), .n31_adj_118(n31_adj_4774), 
            .n30_adj_119(n30_adj_4775), .\d10[70] (d10_adj_5680[70]), .\d10[71] (d10_adj_5680[71]), 
            .n6_adj_120(n6_adj_4831), .n33_adj_121(n33_adj_4772), .n24_adj_122(n24_adj_4804), 
            .n9_adj_123(n9_adj_4828), .n27_adj_124(n27_adj_4801), .n26_adj_125(n26_adj_4802), 
            .n8_adj_126(n8_adj_4829), .n32_adj_127(n32_adj_4773), .n35_adj_128(n35_adj_4770), 
            .n37(n37_adj_4688), .n34_adj_129(n34_adj_4771), .n37_adj_130(n37_adj_4768), 
            .n36(n36_adj_4769), .n29_adj_131(n29_adj_4799), .n19_adj_132(n19_adj_4573), 
            .n28_adj_133(n28_adj_4800), .n31_adj_134(n31_adj_4797), .n30_adj_135(n30_adj_4798), 
            .n33_adj_136(n33_adj_4795), .n36_adj_137(n36_adj_4694), .n118(n118), 
            .n120(n120_adj_5051), .cout(cout_adj_5656), .n32_adj_138(n32_adj_4796), 
            .n35_adj_139(n35_adj_4793), .n34_adj_140(n34_adj_4794), .n37_adj_141(n37_adj_4811), 
            .n18_adj_142(n18_adj_4574), .n36_adj_143(n36_adj_4810), .n115(n115), 
            .n117(n117_adj_5050), .n112(n112), .n114(n114_adj_5049), .\CIC1_outSin[1] (CIC1_outSin[1]), 
            .\CIC1_outSin[2] (CIC1_outSin[2]), .\CIC1_outSin[3] (CIC1_outSin[3]), 
            .\CIC1_outSin[4] (CIC1_outSin[4]), .\CIC1_outSin[5] (CIC1_outSin[5]), 
            .MYLED_0_0(MYLED_0_0), .MYLED_0_1(MYLED_0_1), .MYLED_0_2(MYLED_0_2), 
            .MYLED_0_3(MYLED_0_3), .MYLED_0_4(MYLED_0_4), .MYLED_0_5(MYLED_0_5), 
            .n87_adj_228({n36_adj_5129, n39, n42, n45, n48, n51, 
            n54, n57, n60, n63_adj_5130, n66_adj_5131, n69, n72, 
            n75, n78_adj_5132, n81_adj_5133}), .n29_adj_145(n29_adj_4706), 
            .n109(n109), .n111(n111_adj_5048), .n106(n106), .n108(n108_adj_5047), 
            .n28_adj_146(n28_adj_4707), .n11_adj_147(n11_adj_4826), .n10_adj_148(n10_adj_4827), 
            .n13_adj_149(n13_adj_4824), .n12_adj_150(n12_adj_4825), .n103(n103), 
            .n105(n105_adj_5046), .n3(n3_adj_4763), .n27_adj_151(n27_adj_4708), 
            .n31_adj_152(n31_adj_4704), .n26_adj_153(n26_adj_4709), .n100(n100), 
            .n102(n102_adj_5045), .n2(n2_adj_4764), .n5_adj_154(n5_adj_4761), 
            .n4_adj_155(n4_adj_4762), .n30_adj_156(n30_adj_4705), .n33_adj_157(n33_adj_4702), 
            .n32_adj_158(n32_adj_4703), .n35_adj_159(n35_adj_4700), .n34_adj_160(n34_adj_4701), 
            .n3_adj_161(n3_adj_4568), .n2_adj_162(n2_adj_4569), .n5_adj_163(n5_adj_4730), 
            .n97(n97), .n99(n99_adj_5044), .n4_adj_164(n4_adj_4567), .n63_adj_165(n63), 
            .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_5705[2]), .n7_adj_166(n7_adj_4728), 
            .n6_adj_167(n6_adj_4729), .n9_adj_168(n9_adj_4726), .n8_adj_169(n8_adj_4727), 
            .n11_adj_170(n11_adj_4724), .n10_adj_171(n10_adj_4725), .n64(n64), 
            .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_5705[3]), .n17304(n17304), 
            .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_5705[4]), .n66_adj_172(n66), 
            .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_5705[5]), .n67(n67), 
            .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_5705[6]), .n21_adj_173(n21_adj_4571), 
            .n20_adj_174(n20_adj_4572), .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_5705[7]), 
            .n94(n94), .n96(n96_adj_5043), .n91(n91), .n93(n93_adj_5042), 
            .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_5705[8]), .n23_adj_175(n23_adj_4836), 
            .n22_adj_176(n22_adj_4570), .n88(n88), .n90(n90_adj_5041), 
            .n25_adj_177(n25), .n24_adj_178(n24_adj_4812), .n85(n85), 
            .n87(n87_adj_5040), .n82(n82), .n84(n84_adj_5039), .n79(n79), 
            .n81_adj_179(n81_adj_5038), .n76(n76), .n78_adj_180(n78_adj_5037), 
            .n13_adj_181(n13_adj_4722), .n12_adj_182(n12_adj_4723), .n15_adj_183(n15_adj_4720), 
            .n14_adj_184(n14_adj_4721), .n37_adj_185(n37_adj_4698), .n36_adj_186(n36_adj_4699), 
            .n17_adj_187(n17_adj_4718), .n16_adj_188(n16_adj_4719), .n19_adj_189(n19_adj_4716), 
            .n18_adj_190(n18_adj_4717), .n21_adj_191(n21_adj_4714), .n20_adj_192(n20_adj_4715), 
            .n23_adj_193(n23_adj_4712), .n22_adj_194(n22_adj_4713), .n25_adj_195(n25_adj_4710), 
            .n24_adj_196(n24_adj_4711), .n15_adj_197(n15_adj_4822), .n14_adj_198(n14_adj_4823), 
            .n17_adj_199(n17_adj_4820), .n16_adj_200(n16_adj_4821), .n19_adj_201(n19_adj_4818), 
            .n18_adj_202(n18_adj_4819), .n21_adj_203(n21_adj_4816), .n20_adj_204(n20_adj_4817), 
            .n23_adj_205(n23_adj_4814), .n22_adj_206(n22_adj_4815), .n25_adj_207(n25_adj_4780), 
            .\d10[65] (d10_adj_5680[65]), .\d10[63] (d10_adj_5680[63]), 
            .n3_adj_208(n3_adj_4692), .n2_adj_209(n2_adj_4693), .\d10[64] (d10_adj_5680[64]), 
            .\d10[61] (d10_adj_5680[61]), .\d10[62] (d10_adj_5680[62]), 
            .n17293(n17293), .\d10[59] (d10_adj_5680[59]), .n5_adj_210(n5_adj_4690), 
            .n4_adj_211(n4_adj_4691), .n7_adj_212(n7_adj_4687), .n6_adj_213(n6_adj_4689), 
            .n3_adj_214(n3_adj_4834), .n2_adj_215(n2_adj_4835), .n17317(n17317), 
            .\d10[60] (d10_adj_5680[60]), .n9_adj_216(n9_adj_4655), .n8_adj_217(n8_adj_4658), 
            .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5705[10]), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5705[11]), 
            .n11_adj_218(n11_adj_4617), .n10_adj_219(n10_adj_4625), .n13_adj_220(n13_adj_4579), 
            .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_5705[9]), .n12_adj_221(n12_adj_4592), 
            .n15_adj_222(n15_adj_4577), .n14_adj_223(n14_adj_4578), .n17_adj_224(n17_adj_4575), 
            .n16_adj_225(n16_adj_4576), .n27_adj_226(n27), .n26_adj_227(n26)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(177[45] 183[2])
    CCU2C _add_1_1559_add_4_36 (.A0(d4[69]), .B0(d3[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[70]), .B1(d3[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16055), .COUT(n16056), .S0(n84_adj_5344), .S1(n81_adj_5343));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_3 (.A0(d6[36]), .B0(cout_adj_5341), .C0(n183_adj_4960), 
          .D0(n37_adj_4698), .A1(d6[37]), .B1(cout_adj_5341), .C1(n180_adj_4959), 
          .D1(n36_adj_4699), .CIN(n16002), .COUT(n16003), .S0(d7_71__N_1531[36]), 
          .S1(d7_71__N_1531[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_34 (.A0(d4[67]), .B0(d3[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[68]), .B1(d3[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16054), .COUT(n16055), .S0(n90_adj_5346), .S1(n87_adj_5345));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_34.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i2_rep_174 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(n17750));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(247[8] 297[4])
    defparam o_Rx_Byte_i2_rep_174.GSR = "ENABLED";
    PFUMX i6228 (.BLUT(n17646), .ALUT(n17647), .C0(n17751), .Z(n17648));
    LUT4 mux_325_i25_4_lut (.A(n11959), .B(n247), .C(n17625), .D(n2571), 
         .Z(n2346)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i25_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1559_add_4_32 (.A0(d4[65]), .B0(d3[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[66]), .B1(d3[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16053), .COUT(n16054), .S0(n96_adj_5348), .S1(n93_adj_5347));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_30 (.A0(d4[63]), .B0(d3[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[64]), .B1(d3[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16052), .COUT(n16053), .S0(n102_adj_5350), .S1(n99_adj_5349));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_28 (.A0(d4[61]), .B0(d3[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[62]), .B1(d3[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16051), .COUT(n16052), .S0(n108_adj_5352), .S1(n105_adj_5351));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_26 (.A0(d4[59]), .B0(d3[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[60]), .B1(d3[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16050), .COUT(n16051), .S0(n114_adj_5354), .S1(n111_adj_5353));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5341), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16002));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1463_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1463_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_24 (.A0(d4[57]), .B0(d3[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[58]), .B1(d3[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16049), .COUT(n16050), .S0(n120_adj_5356), .S1(n117_adj_5355));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_24.INJECT1_1 = "NO";
    LUT4 PWMOut_I_0_1_lut (.A(PWMOutP4_c), .Z(PWMOutN4_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(141[19:26])
    defparam PWMOut_I_0_1_lut.init = 16'h5555;
    LUT4 i2272_3_lut_4_lut (.A(n17750), .B(n17630), .C(o_Rx_Byte[3]), 
         .D(n238_adj_5634), .Z(n11961)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam i2272_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1559_add_4_22 (.A0(d4[55]), .B0(d3[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[56]), .B1(d3[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16048), .COUT(n16049), .S0(n126_adj_5358), .S1(n123_adj_5357));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_22.INJECT1_1 = "NO";
    LUT4 mux_325_i26_4_lut (.A(n11961), .B(n244), .C(n17625), .D(n2571), 
         .Z(n2345)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i26_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1559_add_4_20 (.A0(d4[53]), .B0(d3[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[54]), .B1(d3[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16047), .COUT(n16048), .S0(n132_adj_5360), .S1(n129_adj_5359));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_23 (.A0(d6[56]), .B0(cout_adj_5341), .C0(n123_adj_4940), 
          .D0(n17_adj_4718), .A1(d6[57]), .B1(cout_adj_5341), .C1(n120_adj_4939), 
          .D1(n16_adj_4719), .CIN(n16012), .COUT(n16013), .S0(d7_71__N_1531[56]), 
          .S1(d7_71__N_1531[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_18 (.A0(d4[51]), .B0(d3[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[52]), .B1(d3[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16046), .COUT(n16047), .S0(n138_adj_5362), .S1(n135_adj_5361));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_21 (.A0(d6[54]), .B0(cout_adj_5341), .C0(n129_adj_4942), 
          .D0(n19_adj_4716), .A1(d6[55]), .B1(cout_adj_5341), .C1(n126_adj_4941), 
          .D1(n18_adj_4717), .CIN(n16011), .COUT(n16012), .S0(d7_71__N_1531[54]), 
          .S1(d7_71__N_1531[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_16 (.A0(d4[49]), .B0(d3[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[50]), .B1(d3[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16045), .COUT(n16046), .S0(n144_adj_5364), .S1(n141_adj_5363));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_16.INJECT1_1 = "NO";
    SinCos SinCos1 (.clk_80mhz(clk_80mhz), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    CCU2C _add_1_1559_add_4_14 (.A0(d4[47]), .B0(d3[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[48]), .B1(d3[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16044), .COUT(n16045), .S0(n150_adj_5366), .S1(n147_adj_5365));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_12 (.A0(d4[45]), .B0(d3[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[46]), .B1(d3[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16043), .COUT(n16044), .S0(n156_adj_5368), .S1(n153_adj_5367));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_19 (.A0(d6[52]), .B0(cout_adj_5341), .C0(n135_adj_4944), 
          .D0(n21_adj_4714), .A1(d6[53]), .B1(cout_adj_5341), .C1(n132_adj_4943), 
          .D1(n20_adj_4715), .CIN(n16010), .COUT(n16011), .S0(d7_71__N_1531[52]), 
          .S1(d7_71__N_1531[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_10 (.A0(d4[43]), .B0(d3[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[44]), .B1(d3[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16042), .COUT(n16043), .S0(n162_adj_5370), .S1(n159_adj_5369));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_17 (.A0(d6[50]), .B0(cout_adj_5341), .C0(n141_adj_4946), 
          .D0(n23_adj_4712), .A1(d6[51]), .B1(cout_adj_5341), .C1(n138_adj_4945), 
          .D1(n22_adj_4713), .CIN(n16009), .COUT(n16010), .S0(d7_71__N_1531[50]), 
          .S1(d7_71__N_1531[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_8 (.A0(d4[41]), .B0(d3[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[42]), .B1(d3[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16041), .COUT(n16042), .S0(n168_adj_5372), .S1(n165_adj_5371));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_15 (.A0(d6[48]), .B0(cout_adj_5341), .C0(n147_adj_4948), 
          .D0(n25_adj_4710), .A1(d6[49]), .B1(cout_adj_5341), .C1(n144_adj_4947), 
          .D1(n24_adj_4711), .CIN(n16008), .COUT(n16009), .S0(d7_71__N_1531[48]), 
          .S1(d7_71__N_1531[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam _add_1_1463_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_6 (.A0(d4[39]), .B0(d3[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[40]), .B1(d3[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16040), .COUT(n16041), .S0(n174_adj_5374), .S1(n171_adj_5373));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_6.INJECT1_1 = "NO";
    LUT4 mux_325_i23_4_lut (.A(n2548), .B(n253), .C(n17625), .D(n2571), 
         .Z(n2348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i23_4_lut.init = 16'hcfca;
    CCU2C _add_1_1559_add_4_4 (.A0(d4[37]), .B0(d3[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[38]), .B1(d3[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16039), .COUT(n16040), .S0(n180_adj_5376), .S1(n177_adj_5375));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1559_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[36]), .B1(d3[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16039), .S1(n183_adj_5377));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(68[13:20])
    defparam _add_1_1559_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1559_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1559_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_38 (.A0(d_d_tmp[35]), .B0(d_tmp[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16038), .S0(d6_71__N_1459[35]), .S1(cout_adj_5217));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1520_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_38.INJECT1_1 = "NO";
    nco_sig ncoGen (.\phase_accum[63] (phase_accum[63]), .sinGen_c(sinGen_c)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(157[10] 163[2])
    \CIC(width=72,decimation_ratio=4096)_U1  CIC1Cos (.d_tmp({d_tmp_adj_5665}), 
            .clk_80mhz(clk_80mhz), .d5({d5_adj_5671}), .d_d_tmp({d_d_tmp_adj_5666}), 
            .d2({d2_adj_5668}), .d2_71__N_490({d2_71__N_490_adj_5684}), 
            .d3({d3_adj_5669}), .d3_71__N_562({d3_71__N_562_adj_5685}), 
            .d4({d4_adj_5670}), .d4_71__N_634({d4_71__N_634_adj_5686}), 
            .d5_71__N_706({d5_71__N_706_adj_5687}), .d6({d6_adj_5672}), 
            .d6_71__N_1459({d6_71__N_1459_adj_5699}), .d_d6({d_d6_adj_5673}), 
            .d7({d7_adj_5674}), .d7_71__N_1531({d7_71__N_1531_adj_5700}), 
            .d_d7({d_d7_adj_5675}), .d8({d8_adj_5676}), .d8_71__N_1603({d8_71__N_1603_adj_5701}), 
            .d_d8({d_d8_adj_5677}), .d9({d9_adj_5678}), .d9_71__N_1675({d9_71__N_1675_adj_5702}), 
            .d_d9({d_d9_adj_5679}), .CIC1_outCos({CIC1_outCos}), .d1({d1_adj_5667}), 
            .d1_71__N_418({d1_71__N_418_adj_5683}), .count({count_adj_5682}), 
            .n32(n32_adj_4662), .n7(n7), .n6(n6), .\CICGain[1] (CICGain[1]), 
            .\d10[59] (d10_adj_5680[59]), .n17293(n17293), .n33(n33_adj_4584), 
            .n32_adj_1(n32_adj_4585), .\d10[62] (d10_adj_5680[62]), .\d10[63] (d10_adj_5680[63]), 
            .\CICGain[0] (CICGain[0]), .n63(n63), .\d10[60] (d10_adj_5680[60]), 
            .n17317(n17317), .\d10[64] (d10_adj_5680[64]), .n64(n64), 
            .\d10[65] (d10_adj_5680[65]), .n17304(n17304), .\d10[66] (d10_adj_5680[66]), 
            .n66(n66), .n3(n3_adj_4615), .\d10[67] (d10_adj_5680[67]), 
            .n67(n67), .n2(n2_adj_4616), .n35(n35_adj_4582), .n34(n34_adj_4583), 
            .n3_adj_2(n3_adj_2761), .n2_adj_3(n2_adj_2762), .n35_adj_4(n35_adj_4659), 
            .n37(n37_adj_4580), .n36(n36_adj_4581), .\d10[61] (d10_adj_5680[61]), 
            .\d10[68] (d10_adj_5680[68]), .\d10[69] (d10_adj_5680[69]), 
            .\d10[70] (d10_adj_5680[70]), .\d10[71] (d10_adj_5680[71]), 
            .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_5705[2]), .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_5705[3]), 
            .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_5705[4]), .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_5705[5]), 
            .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_5705[6]), .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_5705[7]), 
            .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_5705[8]), .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_5705[9]), 
            .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5705[10]), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5705[11]), 
            .n34_adj_5(n34_adj_4660), .n37_adj_6(n37_adj_4656), .n36_adj_7(n36_adj_4657), 
            .n13(n13_adj_4681), .n12(n12_adj_4685), .n15(n15_adj_4679), 
            .n14(n14_adj_4680), .n17(n17_adj_4677), .n87_adj_114({n36_adj_5138, 
            n39_adj_5139, n42_adj_5140, n45_adj_5141, n48_adj_5142, 
            n51_adj_5143, n54_adj_5144, n57_adj_5145, n60_adj_5146, 
            n63_adj_5147, n66_adj_5148, n69_adj_5149, n72_adj_5150, 
            n75_adj_5151, n78_adj_5152, n81_adj_5153}), .n11(n11_adj_4607), 
            .n5(n5_adj_2759), .n29(n29_adj_4588), .n28(n28_adj_4589), 
            .n4(n4_adj_2760), .n31(n31_adj_4586), .n7_adj_11(n7_adj_2757), 
            .n30(n30_adj_4587), .n6_adj_12(n6_adj_2758), .n9(n9), .n8(n8), 
            .n11_adj_13(n11), .n10(n10), .n13_adj_14(n13), .n12_adj_15(n12), 
            .n15_adj_16(n15), .n14_adj_17(n14), .n9_adj_18(n9_adj_4682), 
            .n17_adj_19(n17), .n16(n16), .n19(n19), .n18(n18), .n118(n118_adj_5535), 
            .n120(n120_adj_4888), .cout(cout_adj_5089), .n115(n115_adj_5534), 
            .n117(n117_adj_4887), .n8_adj_20(n8_adj_4686), .n21(n21), 
            .n16_adj_21(n16_adj_4678), .n19_adj_22(n19_adj_4675), .n10_adj_23(n10_adj_4608), 
            .n18_adj_24(n18_adj_4676), .n21_adj_25(n21_adj_4673), .n15_adj_26(n15_adj_4641), 
            .n20(n20_adj_4674), .n23(n23_adj_4671), .n21_adj_27(n21_adj_4635), 
            .n22(n22_adj_4672), .n20_adj_28(n20_adj_4636), .n23_adj_29(n23_adj_4633), 
            .n22_adj_30(n22_adj_4634), .n25(n25_adj_4631), .n24(n24_adj_4632), 
            .n27(n27_adj_4629), .n26(n26_adj_4630), .n29_adj_31(n29_adj_4627), 
            .n14_adj_32(n14_adj_4642), .n28_adj_33(n28_adj_4628), .n31_adj_34(n31_adj_4624), 
            .n30_adj_35(n30_adj_4626), .n33_adj_36(n33_adj_4622), .n32_adj_37(n32_adj_4623), 
            .n35_adj_38(n35_adj_4620), .n34_adj_39(n34_adj_4621), .n37_adj_40(n37_adj_4618), 
            .n36_adj_41(n36_adj_4619), .n11_adj_42(n11_adj_4684), .n10_adj_43(n10_adj_4683), 
            .n25_adj_44(n25_adj_4669), .n24_adj_45(n24_adj_4670), .n3_adj_46(n3_adj_4653), 
            .n2_adj_47(n2_adj_4654), .n5_adj_48(n5_adj_4651), .n4_adj_49(n4_adj_4652), 
            .n7_adj_50(n7_adj_4649), .n6_adj_51(n6_adj_4650), .n9_adj_52(n9_adj_4647), 
            .n8_adj_53(n8_adj_4648), .n11_adj_54(n11_adj_4645), .n10_adj_55(n10_adj_4646), 
            .n13_adj_56(n13_adj_4643), .n12_adj_57(n12_adj_4644), .n20_adj_58(n20), 
            .n29_adj_59(n29_adj_4665), .n112(n112_adj_5533), .n114(n114_adj_4886), 
            .n23_adj_60(n23), .n22_adj_61(n22), .n28_adj_62(n28_adj_4666), 
            .n25_adj_63(n25_adj_2756), .n31_adj_64(n31_adj_4663), .n24_adj_65(n24), 
            .n109(n109_adj_5532), .n111(n111_adj_4885), .n106(n106_adj_5531), 
            .n108(n108_adj_4884), .n17_adj_66(n17_adj_4639), .n16_adj_67(n16_adj_4640), 
            .n7_adj_68(n7_adj_4611), .n30_adj_69(n30_adj_4664), .n6_adj_70(n6_adj_4612), 
            .n5_adj_71(n5_adj_4613), .n103(n103_adj_5530), .n105(n105_adj_4883), 
            .n19_adj_72(n19_adj_4637), .n4_adj_73(n4_adj_4614), .n27_adj_74(n27_adj_2754), 
            .n100(n100_adj_5529), .n102(n102_adj_4882), .n26_adj_75(n26_adj_2755), 
            .n29_adj_76(n29_adj_2752), .n28_adj_77(n28_adj_2753), .n97(n97_adj_5528), 
            .n99(n99_adj_4881), .n31_adj_78(n31_adj_2750), .n94(n94_adj_5527), 
            .n96(n96_adj_4880), .n91(n91_adj_5526), .n93(n93_adj_4879), 
            .n18_adj_79(n18_adj_4638), .n9_adj_80(n9_adj_4609), .n8_adj_81(n8_adj_4610), 
            .n30_adj_82(n30_adj_2751), .n33_adj_83(n33), .n13_adj_84(n13_adj_4605), 
            .n32_adj_85(n32_adj_2749), .n88(n88_adj_5525), .n90(n90_adj_4878), 
            .n12_adj_86(n12_adj_4606), .n85(n85_adj_5524), .n87(n87_adj_4877), 
            .n35_adj_87(n35), .n34_adj_88(n34), .n82(n82_adj_5523), .n84(n84_adj_4876), 
            .n79(n79_adj_5522), .n81_adj_89(n81_adj_4875), .n76(n76_adj_5521), 
            .n78_adj_90(n78_adj_4874), .n37_adj_91(n37), .n15_adj_92(n15_adj_4603), 
            .n14_adj_93(n14_adj_4604), .n17_adj_94(n17_adj_4601), .n36_adj_95(n36), 
            .n16_adj_96(n16_adj_4602), .n19_adj_97(n19_adj_4599), .n18_adj_98(n18_adj_4600), 
            .n21_adj_99(n21_adj_4597), .n20_adj_100(n20_adj_4598), .n23_adj_101(n23_adj_4595), 
            .n22_adj_102(n22_adj_4596), .n3_adj_103(n3), .n2_adj_104(n2), 
            .n27_adj_105(n27_adj_4667), .n26_adj_106(n26_adj_4668), .n25_adj_107(n25_adj_4593), 
            .n24_adj_108(n24_adj_4594), .n5_adj_109(n5), .n4_adj_110(n4), 
            .n27_adj_111(n27_adj_4590), .n26_adj_112(n26_adj_4591), .n33_adj_113(n33_adj_4661)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(186[45] 192[2])
    CCU2C _add_1_1520_add_4_36 (.A0(d_d_tmp[33]), .B0(d_tmp[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[34]), .B1(d_tmp[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16037), .COUT(n16038), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_34 (.A0(d_d_tmp[31]), .B0(d_tmp[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[32]), .B1(d_tmp[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16036), .COUT(n16037), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_32 (.A0(d_d_tmp[29]), .B0(d_tmp[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[30]), .B1(d_tmp[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16035), .COUT(n16036), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_30 (.A0(d_d_tmp[27]), .B0(d_tmp[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[28]), .B1(d_tmp[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16034), .COUT(n16035), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_37 (.A0(d7_adj_5674[70]), .B0(cout_adj_5254), 
          .C0(n81_adj_5306), .D0(n3_adj_4653), .A1(d7_adj_5674[71]), .B1(cout_adj_5254), 
          .C1(n78_adj_5305), .D1(n2_adj_4654), .CIN(n16209), .S0(d8_71__N_1603_adj_5701[70]), 
          .S1(d8_71__N_1603_adj_5701[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_37.INJECT1_1 = "NO";
    LUT4 mux_325_i24_4_lut (.A(n11957), .B(n250), .C(n17625), .D(n2571), 
         .Z(n2347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(254[2] 296[6])
    defparam mux_325_i24_4_lut.init = 16'hcfca;
    CCU2C _add_1_1520_add_4_28 (.A0(d_d_tmp[25]), .B0(d_tmp[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[26]), .B1(d_tmp[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16033), .COUT(n16034), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_26 (.A0(d_d_tmp[23]), .B0(d_tmp[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[24]), .B1(d_tmp[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16032), .COUT(n16033), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_35 (.A0(d7_adj_5674[68]), .B0(cout_adj_5254), 
          .C0(n87_adj_5308), .D0(n5_adj_4651), .A1(d7_adj_5674[69]), .B1(cout_adj_5254), 
          .C1(n84_adj_5307), .D1(n4_adj_4652), .CIN(n16208), .COUT(n16209), 
          .S0(d8_71__N_1603_adj_5701[68]), .S1(d8_71__N_1603_adj_5701[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_24 (.A0(d_d_tmp[21]), .B0(d_tmp[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[22]), .B1(d_tmp[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16031), .COUT(n16032), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_22 (.A0(d_d_tmp[19]), .B0(d_tmp[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[20]), .B1(d_tmp[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16030), .COUT(n16031), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_33 (.A0(d7_adj_5674[66]), .B0(cout_adj_5254), 
          .C0(n93_adj_5310), .D0(n7_adj_4649), .A1(d7_adj_5674[67]), .B1(cout_adj_5254), 
          .C1(n90_adj_5309), .D1(n6_adj_4650), .CIN(n16207), .COUT(n16208), 
          .S0(d8_71__N_1603_adj_5701[66]), .S1(d8_71__N_1603_adj_5701[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_20 (.A0(d_d_tmp[17]), .B0(d_tmp[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[18]), .B1(d_tmp[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16029), .COUT(n16030), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_20.INJECT1_1 = "NO";
    AMDemodulator AMDemodulator1 (.CIC1_out_clkSin(CIC1_out_clkSin), .\CIC1_outSin[0] (CIC1_outSin[0]), 
            .CIC1_outCos({CIC1_outCos}), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
            .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_0_0(MYLED_0_0), .MYLED_0_1(MYLED_0_1), 
            .MYLED_0_2(MYLED_0_2), .MYLED_0_3(MYLED_0_3), .MYLED_0_4(MYLED_0_4), 
            .MYLED_0_5(MYLED_0_5), .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), 
            .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), 
            .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), 
            .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), 
            .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DemodOut[9] (DemodOut[9]), 
            .\d_out_d_11__N_1876[17] (d_out_d_11__N_1876[17]), .d_out_d_11__N_1875(d_out_d_11__N_1875), 
            .d_out_d_11__N_1879(d_out_d_11__N_1879), .d_out_d_11__N_1877(d_out_d_11__N_1877), 
            .\d_out_d_11__N_1874[17] (d_out_d_11__N_1874[17]), .d_out_d_11__N_1873(d_out_d_11__N_1873), 
            .\ISquare[31] (ISquare[31]), .n209(n209), .\d_out_d_11__N_2335[17] (d_out_d_11__N_2335[17]), 
            .\d_out_d_11__N_2353[17] (d_out_d_11__N_2353[17]), .\d_out_d_11__N_1892[17] (d_out_d_11__N_1892[17]), 
            .\d_out_d_11__N_1890[17] (d_out_d_11__N_1890[17]), .\d_out_d_11__N_1888[17] (d_out_d_11__N_1888[17]), 
            .\d_out_d_11__N_1886[17] (d_out_d_11__N_1886[17]), .\d_out_d_11__N_1884[17] (d_out_d_11__N_1884[17]), 
            .\d_out_d_11__N_1882[17] (d_out_d_11__N_1882[17]), .\d_out_d_11__N_1880[17] (d_out_d_11__N_1880[17]), 
            .\d_out_d_11__N_1878[17] (d_out_d_11__N_1878[17]), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultResult2({MultResult2}), .MultResult1({MultResult1})) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(221[15] 226[10])
    CCU2C _add_1_1520_add_4_18 (.A0(d_d_tmp[15]), .B0(d_tmp[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[16]), .B1(d_tmp[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16028), .COUT(n16029), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_31 (.A0(d7_adj_5674[64]), .B0(cout_adj_5254), 
          .C0(n99_adj_5312), .D0(n9_adj_4647), .A1(d7_adj_5674[65]), .B1(cout_adj_5254), 
          .C1(n96_adj_5311), .D1(n8_adj_4648), .CIN(n16206), .COUT(n16207), 
          .S0(d8_71__N_1603_adj_5701[64]), .S1(d8_71__N_1603_adj_5701[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_31.INJECT1_1 = "NO";
    VLO i1 (.Z(GND_net));
    CCU2C _add_1_1520_add_4_16 (.A0(d_d_tmp[13]), .B0(d_tmp[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[14]), .B1(d_tmp[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16027), .COUT(n16028), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_14 (.A0(d_d_tmp[11]), .B0(d_tmp[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[12]), .B1(d_tmp[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16026), .COUT(n16027), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_29 (.A0(d7_adj_5674[62]), .B0(cout_adj_5254), 
          .C0(n105_adj_5314), .D0(n11_adj_4645), .A1(d7_adj_5674[63]), 
          .B1(cout_adj_5254), .C1(n102_adj_5313), .D1(n10_adj_4646), .CIN(n16205), 
          .COUT(n16206), .S0(d8_71__N_1603_adj_5701[62]), .S1(d8_71__N_1603_adj_5701[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_29.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut_adj_54 (.A(o_Rx_Byte[0]), .B(o_Rx_Byte[6]), 
         .C(n11_adj_4566), .D(MYLED_0_6), .Z(n17098)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(280[4] 294[10])
    defparam i1_3_lut_4_lut_4_lut_adj_54.init = 16'hfff7;
    CCU2C _add_1_1520_add_4_12 (.A0(d_d_tmp[9]), .B0(d_tmp[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[10]), .B1(d_tmp[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16025), .COUT(n16026), .S0(d6_71__N_1459[9]), 
          .S1(d6_71__N_1459[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_10 (.A0(d_d_tmp[7]), .B0(d_tmp[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[8]), .B1(d_tmp[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16024), .COUT(n16025), .S0(d6_71__N_1459[7]), 
          .S1(d6_71__N_1459[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_27 (.A0(d7_adj_5674[60]), .B0(cout_adj_5254), 
          .C0(n111_adj_5316), .D0(n13_adj_4643), .A1(d7_adj_5674[61]), 
          .B1(cout_adj_5254), .C1(n108_adj_5315), .D1(n12_adj_4644), .CIN(n16204), 
          .COUT(n16205), .S0(d8_71__N_1603_adj_5701[60]), .S1(d8_71__N_1603_adj_5701[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam _add_1_1475_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1475_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1475_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1520_add_4_8 (.A0(d_d_tmp[5]), .B0(d_tmp[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[6]), .B1(d_tmp[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16023), .COUT(n16024), .S0(d6_71__N_1459[5]), 
          .S1(d6_71__N_1459[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam _add_1_1520_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1520_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1520_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1520_add_4_8.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (MixerOutSin, clk_80mhz, DiffOut_c, MixerOutCos, RFIn_c, 
            \LOCosine[3] , MixerOutCos_11__N_250, \LOSine[1] , MixerOutSin_11__N_236, 
            \LOCosine[1] , \LOCosine[4] , \LOCosine[5] , \LOCosine[6] , 
            \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , \LOCosine[10] , 
            \LOCosine[11] , \LOCosine[12] , \LOSine[11] , \LOSine[12] , 
            \LOSine[10] , \LOSine[9] , \LOSine[8] , \LOSine[7] , \LOSine[6] , 
            \LOSine[5] , \LOSine[4] , \LOSine[3] , \LOSine[2] , \LOCosine[2] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]MixerOutSin;
    input clk_80mhz;
    output DiffOut_c;
    output [11:0]MixerOutCos;
    input RFIn_c;
    input \LOCosine[3] ;
    input [11:0]MixerOutCos_11__N_250;
    input \LOSine[1] ;
    input [11:0]MixerOutSin_11__N_236;
    input \LOCosine[1] ;
    input \LOCosine[4] ;
    input \LOCosine[5] ;
    input \LOCosine[6] ;
    input \LOCosine[7] ;
    input \LOCosine[8] ;
    input \LOCosine[9] ;
    input \LOCosine[10] ;
    input \LOCosine[11] ;
    input \LOCosine[12] ;
    input \LOSine[11] ;
    input \LOSine[12] ;
    input \LOSine[10] ;
    input \LOSine[9] ;
    input \LOSine[8] ;
    input \LOSine[7] ;
    input \LOSine[6] ;
    input \LOSine[5] ;
    input \LOSine[4] ;
    input \LOSine[3] ;
    input \LOSine[2] ;
    input \LOCosine[2] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    wire [11:0]MixerOutSin_11__N_212;
    
    wire RFInR;
    wire [11:0]MixerOutCos_11__N_224;
    
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_212[0]), .CK(clk_80mhz), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(clk_80mhz), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(23[10] 27[8])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_224[0]), .CK(clk_80mhz), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(clk_80mhz), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(23[10] 27[8])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_212[11]), .CK(clk_80mhz), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_212[10]), .CK(clk_80mhz), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_212[9]), .CK(clk_80mhz), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_212[8]), .CK(clk_80mhz), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_212[7]), .CK(clk_80mhz), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_212[6]), .CK(clk_80mhz), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_212[5]), .CK(clk_80mhz), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_212[4]), .CK(clk_80mhz), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_212[3]), .CK(clk_80mhz), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_212[2]), .CK(clk_80mhz), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_212[1]), .CK(clk_80mhz), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_250[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_236[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_250[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_250[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_250[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_250[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_250[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_250[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_250[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_250[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_250[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_250[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_224[1]), .CK(clk_80mhz), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_236[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_224[2]), .CK(clk_80mhz), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_224[3]), .CK(clk_80mhz), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_224[4]), .CK(clk_80mhz), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_224[5]), .CK(clk_80mhz), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_224[6]), .CK(clk_80mhz), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_224[7]), .CK(clk_80mhz), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_224[8]), .CK(clk_80mhz), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_224[9]), .CK(clk_80mhz), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_224[10]), .CK(clk_80mhz), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_224[11]), .CK(clk_80mhz), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=166, LSE_RLINE=174 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(32[10] 44[8])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_236[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_236[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_236[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_236[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_236[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_236[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_236[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_236[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_236[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_236[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_250[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (\DataInReg[0] , clk_80mhz, \DataInReg_11__N_1856[0] , counter, 
            \DemodOut[9] , \DataInReg[1] , \DataInReg_11__N_1856[1] , 
            \DataInReg[2] , \DataInReg_11__N_1856[2] , \DataInReg[3] , 
            \DataInReg_11__N_1856[3] , \DataInReg[4] , \DataInReg_11__N_1856[4] , 
            \DataInReg[5] , \DataInReg_11__N_1856[5] , \DataInReg[6] , 
            \DataInReg_11__N_1856[6] , \DataInReg[7] , \DataInReg_11__N_1856[7] , 
            \DataInReg[8] , \DataInReg_11__N_1856[8] , \DataInReg[9] , 
            GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output \DataInReg[0] ;
    input clk_80mhz;
    input \DataInReg_11__N_1856[0] ;
    output [9:0]counter;
    input \DemodOut[9] ;
    output \DataInReg[1] ;
    input \DataInReg_11__N_1856[1] ;
    output \DataInReg[2] ;
    input \DataInReg_11__N_1856[2] ;
    output \DataInReg[3] ;
    input \DataInReg_11__N_1856[3] ;
    output \DataInReg[4] ;
    input \DataInReg_11__N_1856[4] ;
    output \DataInReg[5] ;
    input \DataInReg_11__N_1856[5] ;
    output \DataInReg[6] ;
    input \DataInReg_11__N_1856[6] ;
    output \DataInReg[7] ;
    input \DataInReg_11__N_1856[7] ;
    output \DataInReg[8] ;
    input \DataInReg_11__N_1856[8] ;
    output \DataInReg[9] ;
    input GND_net;
    input VCC_net;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    
    wire clk_80mhz_enable_1407;
    wire [9:0]n45;
    wire [11:0]n3954;
    
    wire n12, n17, n15, n11, n16225, n16224, n16223, n16222, 
        n16221;
    
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1856[0] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i1.GSR = "ENABLED";
    FD1S3AX counter_1006__i0 (.D(n45[0]), .CK(clk_80mhz), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i0.GSR = "ENABLED";
    LUT4 i1156_1_lut (.A(\DemodOut[9] ), .Z(n3954[9])) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(26[3] 27[35])
    defparam i1156_1_lut.init = 16'h5555;
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1856[1] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1856[2] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1856[3] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1856[4] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1856[5] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1856[6] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1856[7] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1856[8] ), .SP(clk_80mhz_enable_1407), 
            .CK(clk_80mhz), .Q(\DataInReg[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n3954[9]), .SP(clk_80mhz_enable_1407), .CK(clk_80mhz), 
            .Q(\DataInReg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=195, LSE_RLINE=201 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(23[8] 35[5])
    defparam DataInReg__i10.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[8]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(26[7:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i6174_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(clk_80mhz_enable_1407)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(26[7:19])
    defparam i6174_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(26[7:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(counter[6]), .B(counter[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(26[7:19])
    defparam i5_2_lut.init = 16'heeee;
    FD1S3AX counter_1006__i1 (.D(n45[1]), .CK(clk_80mhz), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i1.GSR = "ENABLED";
    FD1S3AX counter_1006__i2 (.D(n45[2]), .CK(clk_80mhz), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i2.GSR = "ENABLED";
    FD1S3AX counter_1006__i3 (.D(n45[3]), .CK(clk_80mhz), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i3.GSR = "ENABLED";
    FD1S3AX counter_1006__i4 (.D(n45[4]), .CK(clk_80mhz), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i4.GSR = "ENABLED";
    FD1S3AX counter_1006__i5 (.D(n45[5]), .CK(clk_80mhz), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i5.GSR = "ENABLED";
    FD1S3AX counter_1006__i6 (.D(n45[6]), .CK(clk_80mhz), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i6.GSR = "ENABLED";
    FD1S3AX counter_1006__i7 (.D(n45[7]), .CK(clk_80mhz), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i7.GSR = "ENABLED";
    FD1S3AX counter_1006__i8 (.D(n45[8]), .CK(clk_80mhz), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i8.GSR = "ENABLED";
    FD1S3AX counter_1006__i9 (.D(n45[9]), .CK(clk_80mhz), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006__i9.GSR = "ENABLED";
    CCU2C counter_1006_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16225), .S0(n45[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_11.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_11.INIT1 = 16'h0000;
    defparam counter_1006_add_4_11.INJECT1_0 = "NO";
    defparam counter_1006_add_4_11.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16224), .COUT(n16225), .S0(n45[7]), .S1(n45[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_9.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_9.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_9.INJECT1_0 = "NO";
    defparam counter_1006_add_4_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(26[7:19])
    defparam i1_2_lut.init = 16'heeee;
    CCU2C counter_1006_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16223), .COUT(n16224), .S0(n45[5]), .S1(n45[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_7.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_7.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_7.INJECT1_0 = "NO";
    defparam counter_1006_add_4_7.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16222), .COUT(n16223), .S0(n45[3]), .S1(n45[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_5.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_5.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_5.INJECT1_0 = "NO";
    defparam counter_1006_add_4_5.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16221), .COUT(n16222), .S0(n45[1]), .S1(n45[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_3.INIT0 = 16'haaa0;
    defparam counter_1006_add_4_3.INIT1 = 16'haaa0;
    defparam counter_1006_add_4_3.INJECT1_0 = "NO";
    defparam counter_1006_add_4_3.INJECT1_1 = "NO";
    CCU2C counter_1006_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16221), .S1(n45[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/PWM.v(25[14:29])
    defparam counter_1006_add_4_1.INIT0 = 16'h0000;
    defparam counter_1006_add_4_1.INIT1 = 16'h555f;
    defparam counter_1006_add_4_1.INJECT1_0 = "NO";
    defparam counter_1006_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (clk_80mhz, i_Rx_Serial_c, o_Rx_Byte1, 
            o_Rx_DV1, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input clk_80mhz;
    input i_Rx_Serial_c;
    output [7:0]o_Rx_Byte1;
    output o_Rx_DV1;
    input GND_net;
    input VCC_net;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx1/UartClk[2], is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(37[14:21])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    wire [2:0]r_SM_Main;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(43[17:26])
    
    wire n3, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, r_Rx_Data, UartClk_2_enable_17;
    wire [7:0]r_Rx_Byte;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(41[17:26])
    
    wire UartClk_2_enable_2;
    wire [2:0]r_Bit_Index;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(40[17:28])
    
    wire UartClk_2_enable_36, n16921, n1, n13188, n13173, n16778, 
        n17627, n17636, n17619, n13063, n17623, r_Rx_DV_N_2484, 
        n17662, n17624, n17661, n17620, n16827, UartClk_2_enable_9, 
        n17080, n17082, n17074, n17078, UartClk_2_enable_4, UartClk_2_enable_5, 
        n12547, r_Rx_DV_last_N_2483, UartClk_2_enable_6, UartClk_2_enable_7, 
        n16864, UartClk_2_enable_8;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire UartClk_2_enable_10, n17663, n16803;
    wire [15:0]r_Clock_Count;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(39[18:31])
    
    wire n17639, n16477, n20_adj_2748, n17100, UartClk_2_enable_34, 
        n12564, n17090, n17104;
    wire [2:0]n132;
    
    wire n16950, n10, n16971, n13147;
    wire [15:0]n69;
    
    wire n16219, n16218, n16217, n16216, n16215, n16214, n16213, 
        UartClk_2_enable_25, n16212, n16211;
    
    FD1S3IX r_SM_Main_i0 (.D(n3), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(clk_80mhz), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_2), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n16921), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    PFUMX r_SM_Main_2__I_0_69_Mux_0_i3 (.BLUT(n1), .ALUT(n13188), .C0(r_SM_Main[1]), 
          .Z(n3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;
    LUT4 i1_2_lut_rep_158 (.A(n13173), .B(n16778), .Z(n17627)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_158.init = 16'heeee;
    LUT4 i1_2_lut_rep_150_3_lut_4_lut (.A(n13173), .B(n16778), .C(r_SM_Main[0]), 
         .D(n17636), .Z(n17619)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_150_3_lut_4_lut.init = 16'hfff1;
    LUT4 i6168_2_lut_3_lut_4_lut (.A(n13173), .B(n16778), .C(r_SM_Main[0]), 
         .D(n17636), .Z(UartClk_2_enable_17)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i6168_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i3482_3_lut_4_lut (.A(n13173), .B(n16778), .C(r_SM_Main[0]), 
         .D(n13063), .Z(n13188)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i3482_3_lut_4_lut.init = 16'h1e10;
    LUT4 i2341_2_lut_rep_154_3_lut (.A(n13173), .B(n16778), .C(r_SM_Main[0]), 
         .Z(n17623)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i2341_2_lut_rep_154_3_lut.init = 16'hf1f1;
    LUT4 i6116_2_lut_3_lut_4_lut (.A(n13173), .B(n16778), .C(n17636), 
         .D(r_SM_Main[0]), .Z(r_Rx_DV_N_2484)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i6116_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(r_SM_Main[0]), 
         .B(n16778), .C(n13173), .Z(n17662)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h5757;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main[0]), 
         .B(n17624), .C(r_Rx_Data), .Z(n17661)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i6138_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17620), .C(n16827), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_9)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam i6138_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut (.A(n17080), .B(n17082), .C(n17074), .D(n17078), .Z(n16778)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_4_lut.init = 16'hfffe;
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_4), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_5), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2483), .CK(clk_80mhz), .CD(n12547), 
            .Q(o_Rx_DV1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_6), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_7), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    LUT4 i6149_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17620), .C(n16864), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_2)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam i6149_2_lut_3_lut_4_lut.init = 16'h1000;
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_8), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_167 (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .Z(n17636)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_167.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_151_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), 
         .C(n16778), .D(n13173), .Z(n17620)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i1_2_lut_rep_151_3_lut_4_lut.init = 16'hbbbf;
    FD1S3AX UartClk_1007_1031__i0 (.D(n17[0]), .CK(clk_80mhz), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031__i0.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_9), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_10), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i1 (.D(n17663), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(n17627), .CK(UartClk[2]), .CD(n16803), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[4]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[6]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i6079_3_lut_rep_170 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .Z(n17639)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i6079_3_lut_rep_170.init = 16'h8080;
    LUT4 i1_2_lut_rep_155_4_lut (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .D(n16477), .Z(n17624)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_155_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_4_lut (.A(r_Rx_Data), .B(n17639), .C(n16477), .D(r_SM_Main[0]), 
         .Z(n20_adj_2748)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(87[21:38])
    defparam i1_4_lut_4_lut.init = 16'h04ff;
    LUT4 r_SM_Main_2__I_0_69_Mux_0_i1_3_lut_4_lut_4_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), 
         .C(n16477), .D(n17639), .Z(n1)) /* synthesis lut_function=(A (B (C+!(D)))+!A ((C+!(D))+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(87[21:38])
    defparam r_SM_Main_2__I_0_69_Mux_0_i1_3_lut_4_lut_4_lut.init = 16'hd1dd;
    LUT4 i5681_2_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), .Z(n16864)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5681_2_lut.init = 16'h8888;
    LUT4 i6135_2_lut_3_lut_4_lut (.A(r_Bit_Index[0]), .B(n17619), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_10)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(114[17:39])
    defparam i6135_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i6162_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(n17624), 
         .D(n17100), .Z(UartClk_2_enable_34)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam i6162_4_lut.init = 16'h5455;
    LUT4 i1_2_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n17100)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_43 (.A(r_SM_Main[2]), .B(n20_adj_2748), .C(n17627), 
         .D(r_SM_Main[1]), .Z(n12564)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_43.init = 16'h5044;
    LUT4 i6108_4_lut (.A(n17090), .B(n16778), .C(n13173), .D(r_SM_Main[1]), 
         .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i6108_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_44 (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .Z(n17090)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_44.init = 16'heeee;
    LUT4 i1_4_lut_adj_45 (.A(r_Clock_Count[1]), .B(n16778), .C(n17104), 
         .D(r_Clock_Count[6]), .Z(n16477)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_4_lut_adj_45.init = 16'hfffd;
    LUT4 i1_2_lut_adj_46 (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n17104)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_2_lut_adj_46.init = 16'heeee;
    LUT4 i1_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), .C(r_Bit_Index[0]), 
         .Z(n13063)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_47 (.A(n132[2]), .B(n17623), .C(n13063), .D(r_SM_Main[1]), 
         .Z(n16950)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_47.init = 16'h0200;
    LUT4 i1216_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), .C(r_Bit_Index[0]), 
         .Z(n132[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(119[36:54])
    defparam i1216_3_lut.init = 16'h6a6a;
    LUT4 i1_4_lut_adj_48 (.A(n10), .B(n17627), .C(r_SM_Main[0]), .D(r_SM_Main[1]), 
         .Z(n16971)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_48.init = 16'h0800;
    LUT4 i24_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n10)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i24_2_lut.init = 16'h6666;
    LUT4 i6145_2_lut_3_lut_4_lut (.A(r_Bit_Index[0]), .B(n17619), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_5)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(114[17:39])
    defparam i6145_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i6119_3_lut_4_lut (.A(n17627), .B(r_SM_Main[0]), .C(r_Bit_Index[0]), 
         .D(r_SM_Main[1]), .Z(n16921)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam i6119_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_adj_49 (.A(r_Clock_Count[11]), .B(r_Clock_Count[15]), 
         .Z(n17080)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_2_lut_adj_49.init = 16'heeee;
    LUT4 i1_3_lut_adj_50 (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), .C(r_Clock_Count[7]), 
         .Z(n17082)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_3_lut_adj_50.init = 16'hfefe;
    LUT4 i1_2_lut_adj_51 (.A(r_Clock_Count[14]), .B(r_Clock_Count[10]), 
         .Z(n17074)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_2_lut_adj_51.init = 16'heeee;
    LUT4 i6141_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17620), .C(n16827), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_8)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam i6141_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i3469_4_lut (.A(n13147), .B(r_Clock_Count[6]), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[4]), .Z(n13173)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i3469_4_lut.init = 16'hc8c0;
    LUT4 i3443_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n13147)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i3443_3_lut.init = 16'hecec;
    FD1S3AX UartClk_1007_1031__i1 (.D(n17[1]), .CK(clk_80mhz), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031__i1.GSR = "ENABLED";
    FD1S3AX UartClk_1007_1031__i2 (.D(n17[2]), .CK(clk_80mhz), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i0 (.D(n69[0]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i15 (.D(n69[15]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i14 (.D(n69[14]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i14.GSR = "ENABLED";
    CCU2C UartClk_1007_1031_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16219), .S0(n17[1]), .S1(n17[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031_add_4_3.INIT0 = 16'haaa0;
    defparam UartClk_1007_1031_add_4_3.INIT1 = 16'haaa0;
    defparam UartClk_1007_1031_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_1007_1031_add_4_3.INJECT1_1 = "NO";
    CCU2C UartClk_1007_1031_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16219), .S1(n17[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_1007_1031_add_4_1.INIT0 = 16'h0000;
    defparam UartClk_1007_1031_add_4_1.INIT1 = 16'h555f;
    defparam UartClk_1007_1031_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_1007_1031_add_4_1.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16218), .S0(n69[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_17.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_1009_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_17.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16217), .COUT(n16218), .S0(n69[13]), 
          .S1(n69[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_15.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_15.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_15.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_1009__i13 (.D(n69[13]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i13.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_52 (.A(r_Clock_Count[9]), .B(r_Clock_Count[12]), .Z(n17078)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(135[17:47])
    defparam i1_2_lut_adj_52.init = 16'heeee;
    CCU2C r_Clock_Count_1009_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16216), .COUT(n16217), .S0(n69[11]), 
          .S1(n69[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_13.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_13.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_13.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16215), .COUT(n16216), .S0(n69[9]), 
          .S1(n69[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_11.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_11.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_11.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16214), .COUT(n16215), .S0(n69[7]), 
          .S1(n69[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_9.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_9.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_9.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16213), .COUT(n16214), .S0(n69[5]), 
          .S1(n69[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_7.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_7.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_7.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_1009__i12 (.D(n69[12]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i11 (.D(n69[11]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i11.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i10 (.D(n69[10]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i10.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2484), .SP(UartClk_2_enable_25), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    PFUMX i6238 (.BLUT(n17661), .ALUT(n17662), .C0(r_SM_Main[1]), .Z(n17663));
    FD1P3IX r_Clock_Count_1009__i9 (.D(n69[9]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i9.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i8 (.D(n69[8]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i7 (.D(n69[7]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i6 (.D(n69[6]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i6.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i5 (.D(n69[5]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i4 (.D(n69[4]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i3 (.D(n69[3]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i3.GSR = "ENABLED";
    CCU2C r_Clock_Count_1009_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16212), .COUT(n16213), .S0(n69[3]), 
          .S1(n69[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_5.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_5.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_5.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_1009__i2 (.D(n69[2]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i1 (.D(n69[1]), .SP(UartClk_2_enable_34), 
            .CD(n12564), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009__i1.GSR = "ENABLED";
    LUT4 i2840_1_lut (.A(r_Rx_DV), .Z(n12547)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam i2840_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2483)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i6132_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n16803)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i6132_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i6143_2_lut_3_lut_4_lut (.A(r_Bit_Index[0]), .B(n17619), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_6)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(114[17:39])
    defparam i6143_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(n17627), .Z(UartClk_2_enable_25)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;
    defparam i21_4_lut_4_lut.init = 16'h2505;
    LUT4 i6147_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17620), .C(n16864), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_4)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(69[7] 161[14])
    defparam i6147_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i6111_2_lut_3_lut_4_lut (.A(r_Bit_Index[0]), .B(n17619), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_7)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(114[17:39])
    defparam i6111_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_adj_53 (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), .Z(n16827)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_53.init = 16'hbbbb;
    FD1P3AX r_Bit_Index_i2 (.D(n16950), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n16971), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=229, LSE_RLINE=234 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    CCU2C r_Clock_Count_1009_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16211), .COUT(n16212), .S0(n69[1]), 
          .S1(n69[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_3.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_3.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1009_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_3.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1009_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16211), .S1(n69[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_1.INIT0 = 16'h0000;
    defparam r_Clock_Count_1009_add_4_1.INIT1 = 16'h555f;
    defparam r_Clock_Count_1009_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PLL
//

module PLL (osc_clk_c, clk_80mhz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input osc_clk_c;
    output clk_80mhz;
    input GND_net;
    
    wire osc_clk_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(47[13:20])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    
    wire CLKFB_t;
    
    EHXPLLL PLLInst_0 (.CLKI(osc_clk_c), .CLKFB(CLKFB_t), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .PHASELOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .CLKOP(clk_80mhz), .CLKINTFB(CLKFB_t)) /* synthesis FREQUENCY_PIN_CLKOP="83.333333", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="5", LPF_RESISTOR="16", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=127 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(124[5] 127[2])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "INT_OP";
    defparam PLLInst_0.CLKOP_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.PLL_LOCK_DELAY = 200;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.REFIN_RESET = "DISABLED";
    defparam PLLInst_0.SYNC_ENABLE = "DISABLED";
    defparam PLLInst_0.INT_LOCK_STICKY = "ENABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096) 
//

module \CIC(width=72,decimation_ratio=4096)  (d_tmp, clk_80mhz, d5, d_d_tmp, 
            d_d7, n29, n28, d2, d2_71__N_490, d3, d3_71__N_562, 
            n7, d4, d4_71__N_634, d5_71__N_706, d6, d6_71__N_1459, 
            d_d6, CIC1_out_clkSin, d7, d7_71__N_1531, d8, d8_71__N_1603, 
            d_d8, d9, d9_71__N_1675, d_d9, n6, \CIC1_outSin[0] , 
            d1, d1_71__N_418, count, n9, n8, n11, n10, n13, 
            n12, n31, n30, n33, n15, n14, n17, n16, n19, n18, 
            n32, n5, n4, n35, n7_adj_115, n21, n20, n23, n22, 
            n25, n24, n27, n34, \CICGain[1] , \CICGain[0] , \d10[66] , 
            \d10[67] , n26, n29_adj_116, \d10[69] , \d10[68] , n28_adj_117, 
            n31_adj_118, n30_adj_119, \d10[70] , \d10[71] , n6_adj_120, 
            n33_adj_121, n24_adj_122, n9_adj_123, n27_adj_124, n26_adj_125, 
            n8_adj_126, n32_adj_127, n35_adj_128, n37, n34_adj_129, 
            n37_adj_130, n36, n29_adj_131, n19_adj_132, n28_adj_133, 
            n31_adj_134, n30_adj_135, n33_adj_136, n36_adj_137, n118, 
            n120, cout, n32_adj_138, n35_adj_139, n34_adj_140, n37_adj_141, 
            n18_adj_142, n36_adj_143, n115, n117, n112, n114, \CIC1_outSin[1] , 
            \CIC1_outSin[2] , \CIC1_outSin[3] , \CIC1_outSin[4] , \CIC1_outSin[5] , 
            MYLED_0_0, MYLED_0_1, MYLED_0_2, MYLED_0_3, MYLED_0_4, 
            MYLED_0_5, n87_adj_228, n29_adj_145, n109, n111, n106, 
            n108, n28_adj_146, n11_adj_147, n10_adj_148, n13_adj_149, 
            n12_adj_150, n103, n105, n3, n27_adj_151, n31_adj_152, 
            n26_adj_153, n100, n102, n2, n5_adj_154, n4_adj_155, 
            n30_adj_156, n33_adj_157, n32_adj_158, n35_adj_159, n34_adj_160, 
            n3_adj_161, n2_adj_162, n5_adj_163, n97, n99, n4_adj_164, 
            n63_adj_165, \d_out_11__N_1819[2] , n7_adj_166, n6_adj_167, 
            n9_adj_168, n8_adj_169, n11_adj_170, n10_adj_171, n64, 
            \d_out_11__N_1819[3] , n17304, \d_out_11__N_1819[4] , n66_adj_172, 
            \d_out_11__N_1819[5] , n67, \d_out_11__N_1819[6] , n21_adj_173, 
            n20_adj_174, \d_out_11__N_1819[7] , n94, n96, n91, n93, 
            \d_out_11__N_1819[8] , n23_adj_175, n22_adj_176, n88, n90, 
            n25_adj_177, n24_adj_178, n85, n87, n82, n84, n79, 
            n81_adj_179, n76, n78_adj_180, n13_adj_181, n12_adj_182, 
            n15_adj_183, n14_adj_184, n37_adj_185, n36_adj_186, n17_adj_187, 
            n16_adj_188, n19_adj_189, n18_adj_190, n21_adj_191, n20_adj_192, 
            n23_adj_193, n22_adj_194, n25_adj_195, n24_adj_196, n15_adj_197, 
            n14_adj_198, n17_adj_199, n16_adj_200, n19_adj_201, n18_adj_202, 
            n21_adj_203, n20_adj_204, n23_adj_205, n22_adj_206, n25_adj_207, 
            \d10[65] , \d10[63] , n3_adj_208, n2_adj_209, \d10[64] , 
            \d10[61] , \d10[62] , n17293, \d10[59] , n5_adj_210, n4_adj_211, 
            n7_adj_212, n6_adj_213, n3_adj_214, n2_adj_215, n17317, 
            \d10[60] , n9_adj_216, n8_adj_217, \d_out_11__N_1819[10] , 
            \d_out_11__N_1819[11] , n11_adj_218, n10_adj_219, n13_adj_220, 
            \d_out_11__N_1819[9] , n12_adj_221, n15_adj_222, n14_adj_223, 
            n17_adj_224, n16_adj_225, n27_adj_226, n26_adj_227) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d_d7;
    output n29;
    output n28;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output n7;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output CIC1_out_clkSin;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d_d8;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output n6;
    output \CIC1_outSin[0] ;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output [15:0]count;
    output n9;
    output n8;
    output n11;
    output n10;
    output n13;
    output n12;
    output n31;
    output n30;
    output n33;
    output n15;
    output n14;
    output n17;
    output n16;
    output n19;
    output n18;
    output n32;
    output n5;
    output n4;
    output n35;
    output n7_adj_115;
    output n21;
    output n20;
    output n23;
    output n22;
    output n25;
    output n24;
    output n27;
    output n34;
    input \CICGain[1] ;
    input \CICGain[0] ;
    input \d10[66] ;
    input \d10[67] ;
    output n26;
    output n29_adj_116;
    input \d10[69] ;
    input \d10[68] ;
    output n28_adj_117;
    output n31_adj_118;
    output n30_adj_119;
    input \d10[70] ;
    input \d10[71] ;
    output n6_adj_120;
    output n33_adj_121;
    output n24_adj_122;
    output n9_adj_123;
    output n27_adj_124;
    output n26_adj_125;
    output n8_adj_126;
    output n32_adj_127;
    output n35_adj_128;
    output n37;
    output n34_adj_129;
    output n37_adj_130;
    output n36;
    output n29_adj_131;
    output n19_adj_132;
    output n28_adj_133;
    output n31_adj_134;
    output n30_adj_135;
    output n33_adj_136;
    output n36_adj_137;
    input n118;
    input n120;
    input cout;
    output n32_adj_138;
    output n35_adj_139;
    output n34_adj_140;
    output n37_adj_141;
    output n18_adj_142;
    output n36_adj_143;
    input n115;
    input n117;
    input n112;
    input n114;
    output \CIC1_outSin[1] ;
    output \CIC1_outSin[2] ;
    output \CIC1_outSin[3] ;
    output \CIC1_outSin[4] ;
    output \CIC1_outSin[5] ;
    output MYLED_0_0;
    output MYLED_0_1;
    output MYLED_0_2;
    output MYLED_0_3;
    output MYLED_0_4;
    output MYLED_0_5;
    input [15:0]n87_adj_228;
    output n29_adj_145;
    input n109;
    input n111;
    input n106;
    input n108;
    output n28_adj_146;
    output n11_adj_147;
    output n10_adj_148;
    output n13_adj_149;
    output n12_adj_150;
    input n103;
    input n105;
    output n3;
    output n27_adj_151;
    output n31_adj_152;
    output n26_adj_153;
    input n100;
    input n102;
    output n2;
    output n5_adj_154;
    output n4_adj_155;
    output n30_adj_156;
    output n33_adj_157;
    output n32_adj_158;
    output n35_adj_159;
    output n34_adj_160;
    output n3_adj_161;
    output n2_adj_162;
    output n5_adj_163;
    input n97;
    input n99;
    output n4_adj_164;
    input n63_adj_165;
    output \d_out_11__N_1819[2] ;
    output n7_adj_166;
    output n6_adj_167;
    output n9_adj_168;
    output n8_adj_169;
    output n11_adj_170;
    output n10_adj_171;
    input n64;
    output \d_out_11__N_1819[3] ;
    input n17304;
    output \d_out_11__N_1819[4] ;
    input n66_adj_172;
    output \d_out_11__N_1819[5] ;
    input n67;
    output \d_out_11__N_1819[6] ;
    output n21_adj_173;
    output n20_adj_174;
    output \d_out_11__N_1819[7] ;
    input n94;
    input n96;
    input n91;
    input n93;
    output \d_out_11__N_1819[8] ;
    output n23_adj_175;
    output n22_adj_176;
    input n88;
    input n90;
    output n25_adj_177;
    output n24_adj_178;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81_adj_179;
    input n76;
    input n78_adj_180;
    output n13_adj_181;
    output n12_adj_182;
    output n15_adj_183;
    output n14_adj_184;
    output n37_adj_185;
    output n36_adj_186;
    output n17_adj_187;
    output n16_adj_188;
    output n19_adj_189;
    output n18_adj_190;
    output n21_adj_191;
    output n20_adj_192;
    output n23_adj_193;
    output n22_adj_194;
    output n25_adj_195;
    output n24_adj_196;
    output n15_adj_197;
    output n14_adj_198;
    output n17_adj_199;
    output n16_adj_200;
    output n19_adj_201;
    output n18_adj_202;
    output n21_adj_203;
    output n20_adj_204;
    output n23_adj_205;
    output n22_adj_206;
    output n25_adj_207;
    input \d10[65] ;
    input \d10[63] ;
    output n3_adj_208;
    output n2_adj_209;
    input \d10[64] ;
    input \d10[61] ;
    input \d10[62] ;
    input n17293;
    input \d10[59] ;
    output n5_adj_210;
    output n4_adj_211;
    output n7_adj_212;
    output n6_adj_213;
    output n3_adj_214;
    output n2_adj_215;
    input n17317;
    input \d10[60] ;
    output n9_adj_216;
    output n8_adj_217;
    output \d_out_11__N_1819[10] ;
    output \d_out_11__N_1819[11] ;
    output n11_adj_218;
    output n10_adj_219;
    output n13_adj_220;
    output \d_out_11__N_1819[9] ;
    output n12_adj_221;
    output n15_adj_222;
    output n14_adj_223;
    output n17_adj_224;
    output n16_adj_225;
    output n27_adj_226;
    output n26_adj_227;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(86[6:21])
    
    wire clk_80mhz_enable_142, clk_80mhz_enable_65, d_clk_tmp, n12527, 
        v_comb;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    
    wire n17261;
    wire [71:0]d10;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(47[26:29])
    
    wire n17650, n17330, n17649, n17653, n17652, n17148, n16775, 
        n17659, n17319, n17658, n17665, n17664, n17668, n17667, 
        n17671, n17306, n17670, n17311, n17674, n17673, n17677, 
        n17676, n17680, n17679, clk_80mhz_enable_161, d_clk_tmp_N_1831;
    wire [71:0]d10_71__N_1747;
    
    wire n31_adj_2633, n17138, n17142, n17140, clk_80mhz_enable_211, 
        clk_80mhz_enable_261, clk_80mhz_enable_311, clk_80mhz_enable_361, 
        clk_80mhz_enable_411, clk_80mhz_enable_461, clk_80mhz_enable_511, 
        clk_80mhz_enable_561, clk_80mhz_enable_611, clk_80mhz_enable_661, 
        clk_80mhz_enable_711, n12551, n17752, n17269, n17247, n17239, 
        n63_adj_2644, n131, n64_c, n132, n65, n133, n66_adj_2645, 
        n134, n135, n136, n131_adj_2661, n132_adj_2670, n133_adj_2672, 
        n134_adj_2675, n135_adj_2677, n136_adj_2681, n137;
    
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3JX d_clk_tmp_65 (.D(n12527), .CK(clk_80mhz), .PD(clk_80mhz_enable_142), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(clk_80mhz), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_65), 
            .CK(clk_80mhz), .Q(\CIC1_outSin[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_142), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_115)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 i6075_4_lut (.A(count[5]), .B(count[6]), .C(count[2]), .D(count[9]), 
         .Z(n17261)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6075_4_lut.init = 16'h8000;
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    LUT4 i6218_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n17650)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6218_then_3_lut.init = 16'he4e4;
    LUT4 i6218_else_3_lut (.A(n17330), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n17649)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6218_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i210_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[66] ), 
         .C(\d10[67] ), .Z(n17653)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29_adj_116)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i210_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[69] ), 
         .C(\d10[68] ), .Z(n17652)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28_adj_117)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(count[12]), .B(count[11]), .C(n17148), .D(count[15]), 
         .Z(n16775)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17148)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i6206_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n17659)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6206_then_3_lut.init = 16'he4e4;
    LUT4 i6206_else_3_lut (.A(n17319), .B(\CICGain[1] ), .C(d10[59]), 
         .Z(n17658)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6206_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31_adj_118)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30_adj_119)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(\d10[68] ), 
         .C(\d10[70] ), .Z(n17665)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_3_lut (.A(\d10[71] ), .B(\CICGain[1] ), 
         .C(\d10[69] ), .Z(n17664)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_120)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33_adj_121)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(\d10[67] ), .C(\d10[69] ), 
         .Z(n17668)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_122)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_123)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\d10[70] ), .B(\CICGain[1] ), .C(\d10[68] ), 
         .Z(n17667)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_124)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_125)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 i6199_then_3_lut (.A(\CICGain[1] ), .B(d10[67]), .C(d10[65]), 
         .Z(n17671)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6199_then_3_lut.init = 16'he4e4;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_126)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 i6199_else_3_lut (.A(n17306), .B(\CICGain[1] ), .C(d10[66]), 
         .Z(n17670)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6199_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_127)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35_adj_128)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    LUT4 shift_right_31_i212_3_lut_4_lut_then_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[68]), .D(n17311), .Z(n17674)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((D)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_then_4_lut.init = 16'hf791;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[68]), .D(n17311), .Z(n17673)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i212_3_lut_4_lut_else_4_lut.init = 16'he680;
    LUT4 i11_3_lut_4_lut_then_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[67]), .D(n17306), .Z(n17677)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((D)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_then_4_lut.init = 16'hf791;
    LUT4 i11_3_lut_4_lut_else_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[67]), .D(n17306), .Z(n17676)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam i11_3_lut_4_lut_else_4_lut.init = 16'he680;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34_adj_129)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 i6196_then_3_lut (.A(\CICGain[1] ), .B(d10[68]), .C(d10[66]), 
         .Z(n17680)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6196_then_3_lut.init = 16'he4e4;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37_adj_130)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 i6196_else_3_lut (.A(n17311), .B(\CICGain[1] ), .C(d10[67]), 
         .Z(n17679)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6196_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_131)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19_adj_132)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_133)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_134)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30_adj_135)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_136)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_137)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 mux_1251_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i2_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_138)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35_adj_139)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34_adj_140)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_141)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18_adj_142)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_143)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 mux_1251_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i3_3_lut.init = 16'hcaca;
    LUT4 i2820_2_lut (.A(n31_adj_2633), .B(d_clk_tmp), .Z(n12527)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam i2820_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_28 (.A(n17138), .B(n16775), .C(n17142), .D(n17140), 
         .Z(n31_adj_2633)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_28.init = 16'hfffe;
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    LUT4 mux_1251_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i4_3_lut.init = 16'hcaca;
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_161), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_161), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_211), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_261), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_261), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_261), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_311), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_311), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_361), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_361), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_411), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_461), .CK(clk_80mhz), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_461), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_511), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_511), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_561), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_611), .CK(clk_80mhz), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_611), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_661), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_661), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_711), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_711), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\CIC1_outSin[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1819[2]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\CIC1_outSin[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1819[3]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\CIC1_outSin[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1819[4]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\CIC1_outSin[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1819[5]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\CIC1_outSin[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1819[6]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(MYLED_0_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1819[7]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(MYLED_0_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1819[8]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(MYLED_0_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(MYLED_0_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1819[10]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(MYLED_0_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1819[11]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(MYLED_0_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n87_adj_228[2]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_228[3]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_228[4]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_228[5]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_228[6]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_228[7]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_228[8]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_228[9]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_228[10]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(d_clk_tmp_N_1831), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_228[12]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_228[13]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_228[14]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_228[15]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_145)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    FD1S3IX count__i1 (.D(n87_adj_228[1]), .CK(clk_80mhz), .CD(n12551), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17138)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_29 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17142)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_29.init = 16'hfffe;
    LUT4 i1_4_lut_adj_30 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17140)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_30.init = 16'hfffe;
    LUT4 mux_1251_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1251_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i6_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_146)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11_adj_147)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_148)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_149)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_150)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 i6129_2_lut (.A(n31_adj_2633), .B(n17752), .Z(n12551)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam i6129_2_lut.init = 16'hdddd;
    LUT4 i3284_2_lut (.A(n87_adj_228[11]), .B(n31_adj_2633), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(86[13] 89[16])
    defparam i3284_2_lut.init = 16'hbbbb;
    LUT4 i6124_4_lut_rep_176 (.A(n16775), .B(n17269), .C(n17247), .D(n17239), 
         .Z(n17752)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(74[11:40])
    defparam i6124_4_lut_rep_176.init = 16'h4000;
    LUT4 mux_1251_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i7_3_lut.init = 16'hcaca;
    LUT4 i6124_4_lut_rep_177 (.A(n16775), .B(n17269), .C(n17247), .D(n17239), 
         .Z(clk_80mhz_enable_142)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(74[11:40])
    defparam i6124_4_lut_rep_177.init = 16'h4000;
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_2644), .D(n131), .Z(d_out_11__N_1819[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(n132), .Z(d_out_11__N_1819[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(n133), .Z(d_out_11__N_1819[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_2645), .D(n134), .Z(d_out_11__N_1819[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i61_rep_60_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n17330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i61_rep_60_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27_adj_151)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31_adj_152)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_153)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 mux_1251_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i8_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5_adj_154)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4_adj_155)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[66]), .D(n135), .Z(d_out_11__N_1819[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[67]), .D(n136), .Z(d_out_11__N_1819[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30_adj_156)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33_adj_157)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32_adj_158)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_159)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_160)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_161)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_162)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_163)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 mux_1251_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i9_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_164)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_31 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_165), .D(n131_adj_2661), .Z(\d_out_11__N_1819[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_31.init = 16'hfe10;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7_adj_166)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6_adj_167)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_168)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_169)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_170)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_171)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_32 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(n132_adj_2670), .Z(\d_out_11__N_1819[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_32.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_33 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17304), .D(n133_adj_2672), .Z(\d_out_11__N_1819[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_33.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_34 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_172), .D(n134_adj_2675), .Z(\d_out_11__N_1819[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_34.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_35 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(n135_adj_2677), .Z(\d_out_11__N_1819[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_35.init = 16'hfe10;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21_adj_173)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20_adj_174)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_36 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[67] ), .D(n136_adj_2681), .Z(\d_out_11__N_1819[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_36.init = 16'hfe10;
    LUT4 mux_1251_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1251_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i11_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i209_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[68] ), .D(n137), .Z(\d_out_11__N_1819[8] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i209_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_175)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22_adj_176)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 mux_1251_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i12_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25_adj_177)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24_adj_178)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 mux_1251_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1251_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1251_i15_3_lut (.A(n79), .B(n81_adj_179), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1251_i16_3_lut (.A(n76), .B(n78_adj_180), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1251_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13_adj_181)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12_adj_182)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15_adj_183)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14_adj_184)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37_adj_185)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36_adj_186)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17_adj_187)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16_adj_188)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_189)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_190)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_191)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20_adj_192)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23_adj_193)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22_adj_194)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25_adj_195)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24_adj_196)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_2644), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_197)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i62_rep_49_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n17319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i62_rep_49_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17319), .D(d10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 i3222_2_lut (.A(n87_adj_228[0]), .B(n31_adj_2633), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(86[13] 89[16])
    defparam i3222_2_lut.init = 16'hbbbb;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_198)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_199)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_200)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19_adj_201)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_202)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_203)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 i6124_4_lut (.A(n16775), .B(n17269), .C(n17247), .D(n17239), 
         .Z(d_clk_tmp_N_1831)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(74[11:40])
    defparam i6124_4_lut.init = 16'h4000;
    FD1S3AX v_comb_66_rep_181 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_211)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_181.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_191 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_711)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_191.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_180 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_161)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_180.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_190 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_661)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_190.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_189 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_611)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_189.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_188 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_561)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_188.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_204)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23_adj_205)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63_adj_2644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_206)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25_adj_207)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_185 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_411)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_185.GSR = "ENABLED";
    LUT4 shift_right_31_i137_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(\d10[65] ), .Z(n137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut.init = 16'hf960;
    FD1S3AX v_comb_66_rep_186 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_461)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_186.GSR = "ENABLED";
    LUT4 i6083_4_lut (.A(count[0]), .B(n17261), .C(count[4]), .D(count[10]), 
         .Z(n17269)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6083_4_lut.init = 16'h8000;
    FD1S3AX v_comb_66_rep_184 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_361)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_184.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_179 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_65)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_179.GSR = "ENABLED";
    LUT4 shift_right_31_i64_rep_64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i64_rep_64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_37 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17304), .D(\d10[63] ), .Z(n135_adj_2677)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_37.init = 16'hf960;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_208)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_209)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_172), .D(\d10[64] ), .Z(n136_adj_2681)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 i6061_2_lut (.A(count[8]), .B(count[1]), .Z(n17247)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6061_2_lut.init = 16'h8888;
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_38 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_165), .D(\d10[61] ), .Z(n133_adj_2672)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_38.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_39 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(\d10[62] ), .Z(n134_adj_2675)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_39.init = 16'hf960;
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17293), .D(\d10[59] ), .Z(n131_adj_2661)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5_adj_210)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4_adj_211)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7_adj_212)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6_adj_213)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 i6053_2_lut (.A(count[7]), .B(count[3]), .Z(n17239)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6053_2_lut.init = 16'h8888;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3_adj_214)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2_adj_215)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_183 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_311)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_183.GSR = "ENABLED";
    PFUMX i6250 (.BLUT(n17679), .ALUT(n17680), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[9]));
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_182 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_261)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_182.GSR = "ENABLED";
    PFUMX i6248 (.BLUT(n17676), .ALUT(n17677), .C0(d10[70]), .Z(d_out_11__N_1819[10]));
    PFUMX i6246 (.BLUT(n17673), .ALUT(n17674), .C0(d10[71]), .Z(d_out_11__N_1819[11]));
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_40 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17317), .D(\d10[60] ), .Z(n132_adj_2670)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_40.init = 16'hf960;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_216)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_217)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    PFUMX i6244 (.BLUT(n17670), .ALUT(n17671), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[8]));
    PFUMX i6242 (.BLUT(n17667), .ALUT(n17668), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[10] ));
    PFUMX i6240 (.BLUT(n17664), .ALUT(n17665), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[11] ));
    PFUMX i6236 (.BLUT(n17658), .ALUT(n17659), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_218)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10_adj_219)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66_adj_2645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_220)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    PFUMX i6232 (.BLUT(n17652), .ALUT(n17653), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[9] ));
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_221)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15_adj_222)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_41 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17330), .D(d10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_41.init = 16'hf960;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14_adj_223)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_42 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_2645), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_42.init = 16'hf960;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_224)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_225)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    PFUMX i6230 (.BLUT(n17649), .ALUT(n17650), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    LUT4 shift_right_31_i69_rep_36_3_lut (.A(d10[68]), .B(d10[69]), .C(\CICGain[0] ), 
         .Z(n17306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i69_rep_36_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_187 (.D(clk_80mhz_enable_142), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_511)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_187.GSR = "ENABLED";
    LUT4 shift_right_31_i70_rep_41_3_lut (.A(d10[69]), .B(d10[70]), .C(\CICGain[0] ), 
         .Z(n17311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i70_rep_41_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27_adj_226)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26_adj_227)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (clk_80mhz, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_80mhz;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_4_inv, rom_addr0_r_3_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, rom_dout_2_inv, rom_dout_1_inv, co0_1, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_4_inv, rom_dout_3_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_6_inv, rom_dout_5_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_8_inv, rom_dout_7_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_10_inv, rom_dout_9_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_12_inv, rom_dout_11_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_15_inv, 
        rom_dout_14_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_17_inv, 
        rom_dout_16_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_19_inv, 
        rom_dout_18_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_21_inv, 
        rom_dout_20_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_23_inv, 
        rom_dout_22_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_25_inv, 
        rom_dout_24_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    CCU2C neg_rom_addr0_r_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(702[11] 704[71])
    defparam neg_rom_addr0_r_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_0.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
          .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(710[11] 713[42])
    defparam neg_rom_addr0_r_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
          .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(719[11] 722[42])
    defparam neg_rom_addr0_r_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(728[11] 730[73])
    defparam neg_rom_addr0_r_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_3.INJECT1_1 = "NO";
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    CCU2C neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
          .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(874[11] 877[43])
    defparam neg_rom_dout_s_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
          .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(883[11] 886[43])
    defparam neg_rom_dout_s_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_6_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
          .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(892[11] 895[41])
    defparam neg_rom_dout_s_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_8_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
          .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(901[11] 904[41])
    defparam neg_rom_dout_s_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_10_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
          .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(910[11] 913[42])
    defparam neg_rom_dout_s_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_12_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5), .S0(rom_dout_s_n_11), .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(919[11] 922[42])
    defparam neg_rom_dout_s_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_6.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_13_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(936[11] 938[72])
    defparam neg_rom_dout_c_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_0.INJECT1_1 = "NO";
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    CCU2C neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_15_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
          .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(944[11] 947[43])
    defparam neg_rom_dout_c_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_17_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
          .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(953[11] 956[43])
    defparam neg_rom_dout_c_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_19_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
          .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(962[11] 965[43])
    defparam neg_rom_dout_c_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_21_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
          .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(971[11] 974[43])
    defparam neg_rom_dout_c_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_23_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
          .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(980[11] 983[44])
    defparam neg_rom_dout_c_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_25_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5_1), .S0(rom_dout_c_n_11), .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(989[11] 992[44])
    defparam neg_rom_dout_c_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_6.INJECT1_1 = "NO";
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(147[8] 154[2])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    CCU2C neg_rom_dout_s_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=147, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/SinCos.v(866[11] 868[72])
    defparam neg_rom_dout_s_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_0.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module nco_sig
//

module nco_sig (\phase_accum[63] , sinGen_c) /* synthesis syn_module_defined=1 */ ;
    input \phase_accum[63] ;
    output sinGen_c;
    
    
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/NCO.v(32[18:56])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096)_U1 
//

module \CIC(width=72,decimation_ratio=4096)_U1  (d_tmp, clk_80mhz, d5, 
            d_d_tmp, d2, d2_71__N_490, d3, d3_71__N_562, d4, d4_71__N_634, 
            d5_71__N_706, d6, d6_71__N_1459, d_d6, d7, d7_71__N_1531, 
            d_d7, d8, d8_71__N_1603, d_d8, d9, d9_71__N_1675, d_d9, 
            CIC1_outCos, d1, d1_71__N_418, count, n32, n7, n6, 
            \CICGain[1] , \d10[59] , n17293, n33, n32_adj_1, \d10[62] , 
            \d10[63] , \CICGain[0] , n63, \d10[60] , n17317, \d10[64] , 
            n64, \d10[65] , n17304, \d10[66] , n66, n3, \d10[67] , 
            n67, n2, n35, n34, n3_adj_2, n2_adj_3, n35_adj_4, 
            n37, n36, \d10[61] , \d10[68] , \d10[69] , \d10[70] , 
            \d10[71] , \d_out_11__N_1819[2] , \d_out_11__N_1819[3] , \d_out_11__N_1819[4] , 
            \d_out_11__N_1819[5] , \d_out_11__N_1819[6] , \d_out_11__N_1819[7] , 
            \d_out_11__N_1819[8] , \d_out_11__N_1819[9] , \d_out_11__N_1819[10] , 
            \d_out_11__N_1819[11] , n34_adj_5, n37_adj_6, n36_adj_7, 
            n13, n12, n15, n14, n17, n87_adj_114, n11, n5, n29, 
            n28, n4, n31, n7_adj_11, n30, n6_adj_12, n9, n8, 
            n11_adj_13, n10, n13_adj_14, n12_adj_15, n15_adj_16, n14_adj_17, 
            n9_adj_18, n17_adj_19, n16, n19, n18, n118, n120, 
            cout, n115, n117, n8_adj_20, n21, n16_adj_21, n19_adj_22, 
            n10_adj_23, n18_adj_24, n21_adj_25, n15_adj_26, n20, n23, 
            n21_adj_27, n22, n20_adj_28, n23_adj_29, n22_adj_30, n25, 
            n24, n27, n26, n29_adj_31, n14_adj_32, n28_adj_33, n31_adj_34, 
            n30_adj_35, n33_adj_36, n32_adj_37, n35_adj_38, n34_adj_39, 
            n37_adj_40, n36_adj_41, n11_adj_42, n10_adj_43, n25_adj_44, 
            n24_adj_45, n3_adj_46, n2_adj_47, n5_adj_48, n4_adj_49, 
            n7_adj_50, n6_adj_51, n9_adj_52, n8_adj_53, n11_adj_54, 
            n10_adj_55, n13_adj_56, n12_adj_57, n20_adj_58, n29_adj_59, 
            n112, n114, n23_adj_60, n22_adj_61, n28_adj_62, n25_adj_63, 
            n31_adj_64, n24_adj_65, n109, n111, n106, n108, n17_adj_66, 
            n16_adj_67, n7_adj_68, n30_adj_69, n6_adj_70, n5_adj_71, 
            n103, n105, n19_adj_72, n4_adj_73, n27_adj_74, n100, 
            n102, n26_adj_75, n29_adj_76, n28_adj_77, n97, n99, 
            n31_adj_78, n94, n96, n91, n93, n18_adj_79, n9_adj_80, 
            n8_adj_81, n30_adj_82, n33_adj_83, n13_adj_84, n32_adj_85, 
            n88, n90, n12_adj_86, n85, n87, n35_adj_87, n34_adj_88, 
            n82, n84, n79, n81_adj_89, n76, n78_adj_90, n37_adj_91, 
            n15_adj_92, n14_adj_93, n17_adj_94, n36_adj_95, n16_adj_96, 
            n19_adj_97, n18_adj_98, n21_adj_99, n20_adj_100, n23_adj_101, 
            n22_adj_102, n3_adj_103, n2_adj_104, n27_adj_105, n26_adj_106, 
            n25_adj_107, n24_adj_108, n5_adj_109, n4_adj_110, n27_adj_111, 
            n26_adj_112, n33_adj_113) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d_d7;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d_d8;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output [11:0]CIC1_outCos;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output [15:0]count;
    output n32;
    output n7;
    output n6;
    input \CICGain[1] ;
    output \d10[59] ;
    output n17293;
    output n33;
    output n32_adj_1;
    output \d10[62] ;
    output \d10[63] ;
    input \CICGain[0] ;
    output n63;
    output \d10[60] ;
    output n17317;
    output \d10[64] ;
    output n64;
    output \d10[65] ;
    output n17304;
    output \d10[66] ;
    output n66;
    output n3;
    output \d10[67] ;
    output n67;
    output n2;
    output n35;
    output n34;
    output n3_adj_2;
    output n2_adj_3;
    output n35_adj_4;
    output n37;
    output n36;
    output \d10[61] ;
    output \d10[68] ;
    output \d10[69] ;
    output \d10[70] ;
    output \d10[71] ;
    input \d_out_11__N_1819[2] ;
    input \d_out_11__N_1819[3] ;
    input \d_out_11__N_1819[4] ;
    input \d_out_11__N_1819[5] ;
    input \d_out_11__N_1819[6] ;
    input \d_out_11__N_1819[7] ;
    input \d_out_11__N_1819[8] ;
    input \d_out_11__N_1819[9] ;
    input \d_out_11__N_1819[10] ;
    input \d_out_11__N_1819[11] ;
    output n34_adj_5;
    output n37_adj_6;
    output n36_adj_7;
    output n13;
    output n12;
    output n15;
    output n14;
    output n17;
    input [15:0]n87_adj_114;
    output n11;
    output n5;
    output n29;
    output n28;
    output n4;
    output n31;
    output n7_adj_11;
    output n30;
    output n6_adj_12;
    output n9;
    output n8;
    output n11_adj_13;
    output n10;
    output n13_adj_14;
    output n12_adj_15;
    output n15_adj_16;
    output n14_adj_17;
    output n9_adj_18;
    output n17_adj_19;
    output n16;
    output n19;
    output n18;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    output n8_adj_20;
    output n21;
    output n16_adj_21;
    output n19_adj_22;
    output n10_adj_23;
    output n18_adj_24;
    output n21_adj_25;
    output n15_adj_26;
    output n20;
    output n23;
    output n21_adj_27;
    output n22;
    output n20_adj_28;
    output n23_adj_29;
    output n22_adj_30;
    output n25;
    output n24;
    output n27;
    output n26;
    output n29_adj_31;
    output n14_adj_32;
    output n28_adj_33;
    output n31_adj_34;
    output n30_adj_35;
    output n33_adj_36;
    output n32_adj_37;
    output n35_adj_38;
    output n34_adj_39;
    output n37_adj_40;
    output n36_adj_41;
    output n11_adj_42;
    output n10_adj_43;
    output n25_adj_44;
    output n24_adj_45;
    output n3_adj_46;
    output n2_adj_47;
    output n5_adj_48;
    output n4_adj_49;
    output n7_adj_50;
    output n6_adj_51;
    output n9_adj_52;
    output n8_adj_53;
    output n11_adj_54;
    output n10_adj_55;
    output n13_adj_56;
    output n12_adj_57;
    output n20_adj_58;
    output n29_adj_59;
    input n112;
    input n114;
    output n23_adj_60;
    output n22_adj_61;
    output n28_adj_62;
    output n25_adj_63;
    output n31_adj_64;
    output n24_adj_65;
    input n109;
    input n111;
    input n106;
    input n108;
    output n17_adj_66;
    output n16_adj_67;
    output n7_adj_68;
    output n30_adj_69;
    output n6_adj_70;
    output n5_adj_71;
    input n103;
    input n105;
    output n19_adj_72;
    output n4_adj_73;
    output n27_adj_74;
    input n100;
    input n102;
    output n26_adj_75;
    output n29_adj_76;
    output n28_adj_77;
    input n97;
    input n99;
    output n31_adj_78;
    input n94;
    input n96;
    input n91;
    input n93;
    output n18_adj_79;
    output n9_adj_80;
    output n8_adj_81;
    output n30_adj_82;
    output n33_adj_83;
    output n13_adj_84;
    output n32_adj_85;
    input n88;
    input n90;
    output n12_adj_86;
    input n85;
    input n87;
    output n35_adj_87;
    output n34_adj_88;
    input n82;
    input n84;
    input n79;
    input n81_adj_89;
    input n76;
    input n78_adj_90;
    output n37_adj_91;
    output n15_adj_92;
    output n14_adj_93;
    output n17_adj_94;
    output n36_adj_95;
    output n16_adj_96;
    output n19_adj_97;
    output n18_adj_98;
    output n21_adj_99;
    output n20_adj_100;
    output n23_adj_101;
    output n22_adj_102;
    output n3_adj_103;
    output n2_adj_104;
    output n27_adj_105;
    output n26_adj_106;
    output n25_adj_107;
    output n24_adj_108;
    output n5_adj_109;
    output n4_adj_110;
    output n27_adj_111;
    output n26_adj_112;
    output n33_adj_113;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(70[8:17])
    
    wire clk_80mhz_enable_758, clk_80mhz_enable_798, v_comb;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    wire [71:0]d10;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(47[26:29])
    
    wire n17644, n17643, n17656, n17655, count_15__N_1458, clk_80mhz_enable_848, 
        clk_80mhz_enable_898, clk_80mhz_enable_948, clk_80mhz_enable_998, 
        clk_80mhz_enable_1048, clk_80mhz_enable_1098, clk_80mhz_enable_1148, 
        clk_80mhz_enable_1198, clk_80mhz_enable_1248, clk_80mhz_enable_1298, 
        clk_80mhz_enable_1348, clk_80mhz_enable_1398;
    wire [71:0]d10_71__N_1747;
    
    wire n12562, n16769, n17267, n17235, n17227, n31_adj_2517, n17768, 
        n17255, n17174, n17164, n17168, n17166;
    
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_798), 
            .CK(clk_80mhz), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_758), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 i6188_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n17644)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6188_then_3_lut.init = 16'he4e4;
    LUT4 i6188_else_3_lut (.A(n17293), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n17643)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6188_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_1)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 i6183_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n17656)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6183_then_3_lut.init = 16'he4e4;
    LUT4 i6183_else_3_lut (.A(n17317), .B(\CICGain[1] ), .C(\d10[59] ), 
         .Z(n17655)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6183_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i64_3_lut (.A(\d10[63] ), .B(\d10[64] ), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_rep_33_3_lut (.A(\d10[64] ), .B(\d10[65] ), 
         .C(\CICGain[0] ), .Z(n17304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i65_rep_33_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i67_rep_38_3_lut (.A(\d10[66] ), .B(\d10[67] ), 
         .C(\CICGain[0] ), .Z(n67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i67_rep_38_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3_adj_2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2_adj_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_798), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_848), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_848), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_898), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_948), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_948), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_948), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_998), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_998), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_1048), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_1048), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_1048), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_1048), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_1048), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_1048), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_1048), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_1098), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_1148), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_1148), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_1198), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_1198), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_1248), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_1298), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_1298), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_1348), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_1348), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_1398), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_1398), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1819[2] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1819[3] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1819[4] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1819[5] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1819[6] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1819[7] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1819[8] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(\d_out_11__N_1819[9] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1819[10] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1819[11] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37_adj_6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36_adj_7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    FD1S3IX count__i2 (.D(n87_adj_114[2]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_114[3]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_114[4]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_114[5]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_114[6]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_114[7]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_114[8]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_114[9]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_114[10]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(count_15__N_1458), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_114[12]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_114[13]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_114[14]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_114[15]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7_adj_11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6_adj_12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11_adj_13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13_adj_14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12_adj_15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15_adj_16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14_adj_17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17_adj_19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 mux_1250_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i3_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16_adj_21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15_adj_26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21_adj_27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20_adj_28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 i6114_4_lut (.A(n16769), .B(n17267), .C(n17235), .D(n17227), 
         .Z(count_15__N_1458)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(74[11:40])
    defparam i6114_4_lut.init = 16'h4000;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22_adj_30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 i6151_2_lut (.A(n31_adj_2517), .B(n17768), .Z(n12562)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam i6151_2_lut.init = 16'hdddd;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 i3285_2_lut (.A(n87_adj_114[11]), .B(n31_adj_2517), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(86[13] 89[16])
    defparam i3285_2_lut.init = 16'hbbbb;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29_adj_31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14_adj_32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28_adj_33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31_adj_34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33_adj_36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32_adj_37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35_adj_38)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34_adj_39)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37_adj_40)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_41)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_42)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_43)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25_adj_44)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24_adj_45)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_46)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_47)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5_adj_48)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4_adj_49)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7_adj_50)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6_adj_51)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_52)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_53)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_54)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10_adj_55)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_56)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_57)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_200 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1048)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_200.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20_adj_58)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 i6081_4_lut (.A(count[6]), .B(n17255), .C(count[4]), .D(count[10]), 
         .Z(n17267)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6081_4_lut.init = 16'h8000;
    LUT4 i6050_2_lut (.A(count[5]), .B(count[8]), .Z(n17235)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6050_2_lut.init = 16'h8888;
    FD1S3AX v_comb_66_rep_199 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_998)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_199.GSR = "ENABLED";
    LUT4 i6042_2_lut (.A(count[7]), .B(count[3]), .Z(n17227)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6042_2_lut.init = 16'h8888;
    LUT4 i6069_4_lut (.A(count[2]), .B(count[0]), .C(count[1]), .D(count[9]), 
         .Z(n17255)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6069_4_lut.init = 16'h8000;
    FD1S3AX v_comb_66_rep_198 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_948)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_198.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(count[12]), .B(count[11]), .C(n17174), .D(count[15]), 
         .Z(n16769)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    FD1S3AX v_comb_66_rep_197 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_898)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_197.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17174)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3AX v_comb_66_rep_196 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_848)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_196.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_59)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 mux_1250_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i4_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23_adj_60)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22_adj_61)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_62)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_195 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_798)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_195.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_63)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31_adj_64)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_65)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 mux_1250_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i6_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_66)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_67)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_68)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30_adj_69)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_70)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5_adj_71)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 mux_1250_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i7_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19_adj_72)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4_adj_73)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_23_3_lut (.A(\d10[60] ), .B(\d10[61] ), 
         .C(\CICGain[0] ), .Z(n17293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i61_rep_23_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_74)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 mux_1250_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i8_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_75)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_76)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_77)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 i3224_2_lut (.A(n87_adj_114[0]), .B(n31_adj_2517), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(86[13] 89[16])
    defparam i3224_2_lut.init = 16'hbbbb;
    LUT4 mux_1250_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i9_3_lut.init = 16'hcaca;
    LUT4 i6114_4_lut_rep_192 (.A(n16769), .B(n17267), .C(n17235), .D(n17227), 
         .Z(n17768)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(74[11:40])
    defparam i6114_4_lut_rep_192.init = 16'h4000;
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_78)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 mux_1250_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i10_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_25 (.A(n17164), .B(n16769), .C(n17168), .D(n17166), 
         .Z(n31_adj_2517)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_25.init = 16'hfffe;
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17164)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 mux_1250_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i11_3_lut.init = 16'hcaca;
    LUT4 i6114_4_lut_rep_193 (.A(n16769), .B(n17267), .C(n17235), .D(n17227), 
         .Z(clk_80mhz_enable_758)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(74[11:40])
    defparam i6114_4_lut_rep_193.init = 16'h4000;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18_adj_79)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(109[17:26])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_26 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17168)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_26.init = 16'hfffe;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_80)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_81)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30_adj_82)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_27 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17166)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(80[22:52])
    defparam i1_4_lut_adj_27.init = 16'hfffe;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_83)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_84)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_85)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 mux_1250_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i12_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_86)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 mux_1250_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i13_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35_adj_87)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34_adj_88)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 mux_1250_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i15_3_lut (.A(n79), .B(n81_adj_89), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i16_3_lut (.A(n76), .B(n78_adj_90), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(115[18:27])
    defparam mux_1250_i16_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_91)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_92)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_93)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_94)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_95)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(103[17:32])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i62_rep_47_3_lut (.A(\d10[61] ), .B(\d10[62] ), 
         .C(\CICGain[0] ), .Z(n17317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(119[20:47])
    defparam shift_right_31_i62_rep_47_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_96)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19_adj_97)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_98)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_207 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1398)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_207.GSR = "ENABLED";
    PFUMX i6234 (.BLUT(n17655), .ALUT(n17656), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_99)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_206 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1348)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_206.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_100)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23_adj_101)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_102)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_103)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_104)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_205 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1298)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_205.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n87_adj_114[1]), .CK(clk_80mhz), .CD(n12562), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27_adj_105)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_204 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1248)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_204.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_106)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25_adj_107)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24_adj_108)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_109)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_110)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_203 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1198)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_203.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27_adj_111)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    PFUMX i6226 (.BLUT(n17643), .ALUT(n17644), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    FD1S3AX v_comb_66_rep_202 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1148)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_202.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26_adj_112)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(112[17:26])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33_adj_113)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(106[17:26])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_201 (.D(clk_80mhz_enable_758), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1098)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/CIC.v(57[10] 91[8])
    defparam v_comb_66_rep_201.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (CIC1_out_clkSin, \CIC1_outSin[0] , CIC1_outCos, 
            \DataInReg_11__N_1856[0] , \CIC1_outSin[1] , \CIC1_outSin[2] , 
            \CIC1_outSin[3] , \CIC1_outSin[4] , \CIC1_outSin[5] , MYLED_0_0, 
            MYLED_0_1, MYLED_0_2, MYLED_0_3, MYLED_0_4, MYLED_0_5, 
            \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , \DataInReg_11__N_1856[3] , 
            \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , \DataInReg_11__N_1856[6] , 
            \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] , \DemodOut[9] , 
            \d_out_d_11__N_1876[17] , d_out_d_11__N_1875, d_out_d_11__N_1879, 
            d_out_d_11__N_1877, \d_out_d_11__N_1874[17] , d_out_d_11__N_1873, 
            \ISquare[31] , n209, \d_out_d_11__N_2335[17] , \d_out_d_11__N_2353[17] , 
            \d_out_d_11__N_1892[17] , \d_out_d_11__N_1890[17] , \d_out_d_11__N_1888[17] , 
            \d_out_d_11__N_1886[17] , \d_out_d_11__N_1884[17] , \d_out_d_11__N_1882[17] , 
            \d_out_d_11__N_1880[17] , \d_out_d_11__N_1878[17] , VCC_net, 
            GND_net, MultResult2, MultResult1) /* synthesis syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input \CIC1_outSin[0] ;
    input [11:0]CIC1_outCos;
    output \DataInReg_11__N_1856[0] ;
    input \CIC1_outSin[1] ;
    input \CIC1_outSin[2] ;
    input \CIC1_outSin[3] ;
    input \CIC1_outSin[4] ;
    input \CIC1_outSin[5] ;
    input MYLED_0_0;
    input MYLED_0_1;
    input MYLED_0_2;
    input MYLED_0_3;
    input MYLED_0_4;
    input MYLED_0_5;
    output \DataInReg_11__N_1856[1] ;
    output \DataInReg_11__N_1856[2] ;
    output \DataInReg_11__N_1856[3] ;
    output \DataInReg_11__N_1856[4] ;
    output \DataInReg_11__N_1856[5] ;
    output \DataInReg_11__N_1856[6] ;
    output \DataInReg_11__N_1856[7] ;
    output \DataInReg_11__N_1856[8] ;
    output \DemodOut[9] ;
    input \d_out_d_11__N_1876[17] ;
    output d_out_d_11__N_1875;
    output d_out_d_11__N_1879;
    output d_out_d_11__N_1877;
    input \d_out_d_11__N_1874[17] ;
    output d_out_d_11__N_1873;
    input \ISquare[31] ;
    output n209;
    input \d_out_d_11__N_2335[17] ;
    input \d_out_d_11__N_2353[17] ;
    input \d_out_d_11__N_1892[17] ;
    input \d_out_d_11__N_1890[17] ;
    input \d_out_d_11__N_1888[17] ;
    input \d_out_d_11__N_1886[17] ;
    input \d_out_d_11__N_1884[17] ;
    input \d_out_d_11__N_1882[17] ;
    input \d_out_d_11__N_1880[17] ;
    input \d_out_d_11__N_1878[17] ;
    input VCC_net;
    input GND_net;
    output [23:0]MultResult2;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(86[6:21])
    wire [11:0]MultDataB;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(29[21:30])
    wire [11:0]MultDataC;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(33[21:30])
    wire [15:0]d_out_d;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(20[21:28])
    wire [17:0]d_out_d_11__N_1894;
    
    wire d_out_d_11__N_1891, d_out_d_11__N_1889, d_out_d_11__N_1887, d_out_d_11__N_1885, 
        d_out_d_11__N_1883, d_out_d_11__N_1881;
    
    FD1S3AX MultDataB_i0 (.D(\CIC1_outSin[0] ), .CK(CIC1_out_clkSin), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i0.GSR = "ENABLED";
    FD1S3AX MultDataC_i0 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), .Q(MultDataC[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i0.GSR = "ENABLED";
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i1.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    FD1S3AX MultDataB_i1 (.D(\CIC1_outSin[1] ), .CK(CIC1_out_clkSin), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i1.GSR = "ENABLED";
    FD1S3AX MultDataB_i2 (.D(\CIC1_outSin[2] ), .CK(CIC1_out_clkSin), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i2.GSR = "ENABLED";
    FD1S3AX MultDataB_i3 (.D(\CIC1_outSin[3] ), .CK(CIC1_out_clkSin), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i3.GSR = "ENABLED";
    FD1S3AX MultDataB_i4 (.D(\CIC1_outSin[4] ), .CK(CIC1_out_clkSin), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i4.GSR = "ENABLED";
    FD1S3AX MultDataB_i5 (.D(\CIC1_outSin[5] ), .CK(CIC1_out_clkSin), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i5.GSR = "ENABLED";
    FD1S3AX MultDataB_i6 (.D(MYLED_0_0), .CK(CIC1_out_clkSin), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i6.GSR = "ENABLED";
    FD1S3AX MultDataB_i7 (.D(MYLED_0_1), .CK(CIC1_out_clkSin), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i7.GSR = "ENABLED";
    FD1S3AX MultDataB_i8 (.D(MYLED_0_2), .CK(CIC1_out_clkSin), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i8.GSR = "ENABLED";
    FD1S3AX MultDataB_i9 (.D(MYLED_0_3), .CK(CIC1_out_clkSin), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i9.GSR = "ENABLED";
    FD1S3AX MultDataB_i10 (.D(MYLED_0_4), .CK(CIC1_out_clkSin), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i10.GSR = "ENABLED";
    FD1S3AX MultDataB_i11 (.D(MYLED_0_5), .CK(CIC1_out_clkSin), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataB_i11.GSR = "ENABLED";
    FD1S3AX MultDataC_i1 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), .Q(MultDataC[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i1.GSR = "ENABLED";
    FD1S3AX MultDataC_i2 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), .Q(MultDataC[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i2.GSR = "ENABLED";
    FD1S3AX MultDataC_i3 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), .Q(MultDataC[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i3.GSR = "ENABLED";
    FD1S3AX MultDataC_i4 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), .Q(MultDataC[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i4.GSR = "ENABLED";
    FD1S3AX MultDataC_i5 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), .Q(MultDataC[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i5.GSR = "ENABLED";
    FD1S3AX MultDataC_i6 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), .Q(MultDataC[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i6.GSR = "ENABLED";
    FD1S3AX MultDataC_i7 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), .Q(MultDataC[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i7.GSR = "ENABLED";
    FD1S3AX MultDataC_i8 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), .Q(MultDataC[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i8.GSR = "ENABLED";
    FD1S3AX MultDataC_i9 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), .Q(MultDataC[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i9.GSR = "ENABLED";
    FD1S3AX MultDataC_i10 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), .Q(MultDataC[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i10.GSR = "ENABLED";
    FD1S3AX MultDataC_i11 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), .Q(MultDataC[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam MultDataC_i11.GSR = "ENABLED";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=221, LSE_RLINE=226 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_i10.GSR = "ENABLED";
    LUT4 d_out_d_11__I_2_1_lut (.A(\d_out_d_11__N_1876[17] ), .Z(d_out_d_11__N_1875)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1891), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1889), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1887), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1885), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1883), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1881), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1879), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1877), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1875), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(86[9] 95[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    LUT4 d_out_d_11__I_1_1_lut (.A(\d_out_d_11__N_1874[17] ), .Z(d_out_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    LUT4 i1339_1_lut (.A(\ISquare[31] ), .Z(n209)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1339_1_lut.init = 16'h5555;
    LUT4 mux_81_i1_3_lut (.A(\d_out_d_11__N_2335[17] ), .B(\d_out_d_11__N_2353[17] ), 
         .C(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1894[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(60[11:28])
    defparam mux_81_i1_3_lut.init = 16'h3535;
    LUT4 d_out_d_11__I_10_1_lut (.A(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1891)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_9_1_lut (.A(\d_out_d_11__N_1890[17] ), .Z(d_out_d_11__N_1889)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(\d_out_d_11__N_1888[17] ), .Z(d_out_d_11__N_1887)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(\d_out_d_11__N_1886[17] ), .Z(d_out_d_11__N_1885)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(\d_out_d_11__N_1884[17] ), .Z(d_out_d_11__N_1883)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(\d_out_d_11__N_1882[17] ), .Z(d_out_d_11__N_1881)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_4_1_lut (.A(\d_out_d_11__N_1880[17] ), .Z(d_out_d_11__N_1879)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(\d_out_d_11__N_1878[17] ), .Z(d_out_d_11__N_1877)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(61[22:28])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    Multiplier Multiplier2 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataC({MultDataC}), .MultResult2({MultResult2})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(77[14] 83[27])
    Multiplier_U0 Multiplier1 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataB({MultDataB}), .MultResult1({MultResult1})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/AMDemod.v(69[14] 75[27])
    
endmodule
//
// Verilog Description of module Multiplier
//

module Multiplier (CIC1_out_clkSin, VCC_net, GND_net, MultDataC, MultResult2) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataC;
    output [23:0]MultResult2;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(86[6:21])
    
    MULT18X18D dsp_mult_0 (.A17(MultDataC[11]), .A16(MultDataC[10]), .A15(MultDataC[9]), 
            .A14(MultDataC[8]), .A13(MultDataC[7]), .A12(MultDataC[6]), 
            .A11(MultDataC[5]), .A10(MultDataC[4]), .A9(MultDataC[3]), 
            .A8(MultDataC[2]), .A7(MultDataC[1]), .A6(MultDataC[0]), .A5(GND_net), 
            .A4(GND_net), .A3(GND_net), .A2(GND_net), .A1(GND_net), 
            .A0(GND_net), .B17(MultDataC[11]), .B16(MultDataC[10]), .B15(MultDataC[9]), 
            .B14(MultDataC[8]), .B13(MultDataC[7]), .B12(MultDataC[6]), 
            .B11(MultDataC[5]), .B10(MultDataC[4]), .B9(MultDataC[3]), 
            .B8(MultDataC[2]), .B7(MultDataC[1]), .B6(MultDataC[0]), .B5(GND_net), 
            .B4(GND_net), .B3(GND_net), .B2(GND_net), .B1(GND_net), 
            .B0(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(CIC1_out_clkSin), .CE3(VCC_net), 
            .CE2(VCC_net), .CE1(VCC_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .P35(MultResult2[23]), 
            .P34(MultResult2[22]), .P33(MultResult2[21]), .P32(MultResult2[20]), 
            .P31(MultResult2[19]), .P30(MultResult2[18]), .P29(MultResult2[17]), 
            .P28(MultResult2[16]), .P27(MultResult2[15]), .P26(MultResult2[14]), 
            .P25(MultResult2[13]), .P24(MultResult2[12]), .P23(MultResult2[11]), 
            .P22(MultResult2[10]), .P21(MultResult2[9]), .P20(MultResult2[8]), 
            .P19(MultResult2[7]), .P18(MultResult2[6]), .P17(MultResult2[5]), 
            .P16(MultResult2[4]), .P15(MultResult2[3]), .P14(MultResult2[2]), 
            .P13(MultResult2[1]), .P12(MultResult2[0])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Multiplier.v(84[16] 140[57])
    defparam dsp_mult_0.REG_INPUTA_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTA_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTA_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTB_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTB_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTB_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTC_CLK = "NONE";
    defparam dsp_mult_0.REG_INPUTC_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTC_RST = "RST0";
    defparam dsp_mult_0.REG_PIPELINE_CLK = "CLK0";
    defparam dsp_mult_0.REG_PIPELINE_CE = "CE0";
    defparam dsp_mult_0.REG_PIPELINE_RST = "RST0";
    defparam dsp_mult_0.REG_OUTPUT_CLK = "CLK0";
    defparam dsp_mult_0.REG_OUTPUT_CE = "CE0";
    defparam dsp_mult_0.REG_OUTPUT_RST = "RST0";
    defparam dsp_mult_0.CLK0_DIV = "ENABLED";
    defparam dsp_mult_0.CLK1_DIV = "ENABLED";
    defparam dsp_mult_0.CLK2_DIV = "ENABLED";
    defparam dsp_mult_0.CLK3_DIV = "ENABLED";
    defparam dsp_mult_0.HIGHSPEED_CLK = "NONE";
    defparam dsp_mult_0.GSR = "ENABLED";
    defparam dsp_mult_0.CAS_MATCH_REG = "FALSE";
    defparam dsp_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam dsp_mult_0.MULT_BYPASS = "DISABLED";
    defparam dsp_mult_0.RESETMODE = "ASYNC";
    
endmodule
//
// Verilog Description of module Multiplier_U0
//

module Multiplier_U0 (CIC1_out_clkSin, VCC_net, GND_net, MultDataB, 
            MultResult1) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/top.v(86[6:21])
    
    MULT18X18D dsp_mult_0 (.A17(MultDataB[11]), .A16(MultDataB[10]), .A15(MultDataB[9]), 
            .A14(MultDataB[8]), .A13(MultDataB[7]), .A12(MultDataB[6]), 
            .A11(MultDataB[5]), .A10(MultDataB[4]), .A9(MultDataB[3]), 
            .A8(MultDataB[2]), .A7(MultDataB[1]), .A6(MultDataB[0]), .A5(GND_net), 
            .A4(GND_net), .A3(GND_net), .A2(GND_net), .A1(GND_net), 
            .A0(GND_net), .B17(MultDataB[11]), .B16(MultDataB[10]), .B15(MultDataB[9]), 
            .B14(MultDataB[8]), .B13(MultDataB[7]), .B12(MultDataB[6]), 
            .B11(MultDataB[5]), .B10(MultDataB[4]), .B9(MultDataB[3]), 
            .B8(MultDataB[2]), .B7(MultDataB[1]), .B6(MultDataB[0]), .B5(GND_net), 
            .B4(GND_net), .B3(GND_net), .B2(GND_net), .B1(GND_net), 
            .B0(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(CIC1_out_clkSin), .CE3(VCC_net), 
            .CE2(VCC_net), .CE1(VCC_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .P35(MultResult1[23]), 
            .P34(MultResult1[22]), .P33(MultResult1[21]), .P32(MultResult1[20]), 
            .P31(MultResult1[19]), .P30(MultResult1[18]), .P29(MultResult1[17]), 
            .P28(MultResult1[16]), .P27(MultResult1[15]), .P26(MultResult1[14]), 
            .P25(MultResult1[13]), .P24(MultResult1[12]), .P23(MultResult1[11]), 
            .P22(MultResult1[10]), .P21(MultResult1[9]), .P20(MultResult1[8]), 
            .P19(MultResult1[7]), .P18(MultResult1[6]), .P17(MultResult1[5]), 
            .P16(MultResult1[4]), .P15(MultResult1[3]), .P14(MultResult1[2]), 
            .P13(MultResult1[1]), .P12(MultResult1[0])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/OriginalVersion/impl1/source/Multiplier.v(84[16] 140[57])
    defparam dsp_mult_0.REG_INPUTA_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTA_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTA_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTB_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTB_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTB_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTC_CLK = "NONE";
    defparam dsp_mult_0.REG_INPUTC_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTC_RST = "RST0";
    defparam dsp_mult_0.REG_PIPELINE_CLK = "CLK0";
    defparam dsp_mult_0.REG_PIPELINE_CE = "CE0";
    defparam dsp_mult_0.REG_PIPELINE_RST = "RST0";
    defparam dsp_mult_0.REG_OUTPUT_CLK = "CLK0";
    defparam dsp_mult_0.REG_OUTPUT_CE = "CE0";
    defparam dsp_mult_0.REG_OUTPUT_RST = "RST0";
    defparam dsp_mult_0.CLK0_DIV = "ENABLED";
    defparam dsp_mult_0.CLK1_DIV = "ENABLED";
    defparam dsp_mult_0.CLK2_DIV = "ENABLED";
    defparam dsp_mult_0.CLK3_DIV = "ENABLED";
    defparam dsp_mult_0.HIGHSPEED_CLK = "NONE";
    defparam dsp_mult_0.GSR = "ENABLED";
    defparam dsp_mult_0.CAS_MATCH_REG = "FALSE";
    defparam dsp_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam dsp_mult_0.MULT_BYPASS = "DISABLED";
    defparam dsp_mult_0.RESETMODE = "ASYNC";
    
endmodule
