module simpleSine(
    clk,
    rst,
    sample_clock_ce,
    phase_inc_carrGen,
    sinewave
);


parameter SB = 12, // SINE_BITS
          PB = 64; // PHASE_BITS

input clk;
input wire rst;
input wire sample_clock_ce;
input reg signed [PB-1:0] phase_inc_carrGen;
output reg signed[SB-1:0] sinewave;

reg [PB-1:0] phase = 0;

always @(posedge clk or posedge rst) begin
    if (rst)
        phase <= 0;
    else if (sample_clock_ce)
        phase <= phase + phase_inc_carrGen;
end

always @(posedge clk) begin
	if (sample_clock_ce) begin
        case(phase[63:52])
        12'h000: sinewave <= 12'h000;
        12'h001: sinewave <= 12'h003;
        12'h002: sinewave <= 12'h006;
        12'h003: sinewave <= 12'h009;
        12'h004: sinewave <= 12'h00C;
        12'h005: sinewave <= 12'h00F;
        12'h006: sinewave <= 12'h012;
        12'h007: sinewave <= 12'h015;
        12'h008: sinewave <= 12'h019;
        12'h009: sinewave <= 12'h01C;
        12'h00A: sinewave <= 12'h01F;
        12'h00B: sinewave <= 12'h022;
        12'h00C: sinewave <= 12'h025;
        12'h00D: sinewave <= 12'h028;
        12'h00E: sinewave <= 12'h02B;
        12'h00F: sinewave <= 12'h02F;
        12'h010: sinewave <= 12'h032;
        12'h011: sinewave <= 12'h035;
        12'h012: sinewave <= 12'h038;
        12'h013: sinewave <= 12'h03B;
        12'h014: sinewave <= 12'h03E;
        12'h015: sinewave <= 12'h041;
        12'h016: sinewave <= 12'h045;
        12'h017: sinewave <= 12'h048;
        12'h018: sinewave <= 12'h04B;
        12'h019: sinewave <= 12'h04E;
        12'h01A: sinewave <= 12'h051;
        12'h01B: sinewave <= 12'h054;
        12'h01C: sinewave <= 12'h057;
        12'h01D: sinewave <= 12'h05B;
        12'h01E: sinewave <= 12'h05E;
        12'h01F: sinewave <= 12'h061;
        12'h020: sinewave <= 12'h064;
        12'h021: sinewave <= 12'h067;
        12'h022: sinewave <= 12'h06A;
        12'h023: sinewave <= 12'h06D;
        12'h024: sinewave <= 12'h070;
        12'h025: sinewave <= 12'h074;
        12'h026: sinewave <= 12'h077;
        12'h027: sinewave <= 12'h07A;
        12'h028: sinewave <= 12'h07D;
        12'h029: sinewave <= 12'h080;
        12'h02A: sinewave <= 12'h083;
        12'h02B: sinewave <= 12'h086;
        12'h02C: sinewave <= 12'h08A;
        12'h02D: sinewave <= 12'h08D;
        12'h02E: sinewave <= 12'h090;
        12'h02F: sinewave <= 12'h093;
        12'h030: sinewave <= 12'h096;
        12'h031: sinewave <= 12'h099;
        12'h032: sinewave <= 12'h09C;
        12'h033: sinewave <= 12'h09F;
        12'h034: sinewave <= 12'h0A3;
        12'h035: sinewave <= 12'h0A6;
        12'h036: sinewave <= 12'h0A9;
        12'h037: sinewave <= 12'h0AC;
        12'h038: sinewave <= 12'h0AF;
        12'h039: sinewave <= 12'h0B2;
        12'h03A: sinewave <= 12'h0B5;
        12'h03B: sinewave <= 12'h0B9;
        12'h03C: sinewave <= 12'h0BC;
        12'h03D: sinewave <= 12'h0BF;
        12'h03E: sinewave <= 12'h0C2;
        12'h03F: sinewave <= 12'h0C5;
        12'h040: sinewave <= 12'h0C8;
        12'h041: sinewave <= 12'h0CB;
        12'h042: sinewave <= 12'h0CE;
        12'h043: sinewave <= 12'h0D2;
        12'h044: sinewave <= 12'h0D5;
        12'h045: sinewave <= 12'h0D8;
        12'h046: sinewave <= 12'h0DB;
        12'h047: sinewave <= 12'h0DE;
        12'h048: sinewave <= 12'h0E1;
        12'h049: sinewave <= 12'h0E4;
        12'h04A: sinewave <= 12'h0E7;
        12'h04B: sinewave <= 12'h0EA;
        12'h04C: sinewave <= 12'h0EE;
        12'h04D: sinewave <= 12'h0F1;
        12'h04E: sinewave <= 12'h0F4;
        12'h04F: sinewave <= 12'h0F7;
        12'h050: sinewave <= 12'h0FA;
        12'h051: sinewave <= 12'h0FD;
        12'h052: sinewave <= 12'h100;
        12'h053: sinewave <= 12'h103;
        12'h054: sinewave <= 12'h107;
        12'h055: sinewave <= 12'h10A;
        12'h056: sinewave <= 12'h10D;
        12'h057: sinewave <= 12'h110;
        12'h058: sinewave <= 12'h113;
        12'h059: sinewave <= 12'h116;
        12'h05A: sinewave <= 12'h119;
        12'h05B: sinewave <= 12'h11C;
        12'h05C: sinewave <= 12'h11F;
        12'h05D: sinewave <= 12'h123;
        12'h05E: sinewave <= 12'h126;
        12'h05F: sinewave <= 12'h129;
        12'h060: sinewave <= 12'h12C;
        12'h061: sinewave <= 12'h12F;
        12'h062: sinewave <= 12'h132;
        12'h063: sinewave <= 12'h135;
        12'h064: sinewave <= 12'h138;
        12'h065: sinewave <= 12'h13B;
        12'h066: sinewave <= 12'h13E;
        12'h067: sinewave <= 12'h142;
        12'h068: sinewave <= 12'h145;
        12'h069: sinewave <= 12'h148;
        12'h06A: sinewave <= 12'h14B;
        12'h06B: sinewave <= 12'h14E;
        12'h06C: sinewave <= 12'h151;
        12'h06D: sinewave <= 12'h154;
        12'h06E: sinewave <= 12'h157;
        12'h06F: sinewave <= 12'h15A;
        12'h070: sinewave <= 12'h15D;
        12'h071: sinewave <= 12'h161;
        12'h072: sinewave <= 12'h164;
        12'h073: sinewave <= 12'h167;
        12'h074: sinewave <= 12'h16A;
        12'h075: sinewave <= 12'h16D;
        12'h076: sinewave <= 12'h170;
        12'h077: sinewave <= 12'h173;
        12'h078: sinewave <= 12'h176;
        12'h079: sinewave <= 12'h179;
        12'h07A: sinewave <= 12'h17C;
        12'h07B: sinewave <= 12'h17F;
        12'h07C: sinewave <= 12'h183;
        12'h07D: sinewave <= 12'h186;
        12'h07E: sinewave <= 12'h189;
        12'h07F: sinewave <= 12'h18C;
        12'h080: sinewave <= 12'h18F;
        12'h081: sinewave <= 12'h192;
        12'h082: sinewave <= 12'h195;
        12'h083: sinewave <= 12'h198;
        12'h084: sinewave <= 12'h19B;
        12'h085: sinewave <= 12'h19E;
        12'h086: sinewave <= 12'h1A1;
        12'h087: sinewave <= 12'h1A4;
        12'h088: sinewave <= 12'h1A7;
        12'h089: sinewave <= 12'h1AB;
        12'h08A: sinewave <= 12'h1AE;
        12'h08B: sinewave <= 12'h1B1;
        12'h08C: sinewave <= 12'h1B4;
        12'h08D: sinewave <= 12'h1B7;
        12'h08E: sinewave <= 12'h1BA;
        12'h08F: sinewave <= 12'h1BD;
        12'h090: sinewave <= 12'h1C0;
        12'h091: sinewave <= 12'h1C3;
        12'h092: sinewave <= 12'h1C6;
        12'h093: sinewave <= 12'h1C9;
        12'h094: sinewave <= 12'h1CC;
        12'h095: sinewave <= 12'h1CF;
        12'h096: sinewave <= 12'h1D2;
        12'h097: sinewave <= 12'h1D5;
        12'h098: sinewave <= 12'h1D8;
        12'h099: sinewave <= 12'h1DC;
        12'h09A: sinewave <= 12'h1DF;
        12'h09B: sinewave <= 12'h1E2;
        12'h09C: sinewave <= 12'h1E5;
        12'h09D: sinewave <= 12'h1E8;
        12'h09E: sinewave <= 12'h1EB;
        12'h09F: sinewave <= 12'h1EE;
        12'h0A0: sinewave <= 12'h1F1;
        12'h0A1: sinewave <= 12'h1F4;
        12'h0A2: sinewave <= 12'h1F7;
        12'h0A3: sinewave <= 12'h1FA;
        12'h0A4: sinewave <= 12'h1FD;
        12'h0A5: sinewave <= 12'h200;
        12'h0A6: sinewave <= 12'h203;
        12'h0A7: sinewave <= 12'h206;
        12'h0A8: sinewave <= 12'h209;
        12'h0A9: sinewave <= 12'h20C;
        12'h0AA: sinewave <= 12'h20F;
        12'h0AB: sinewave <= 12'h212;
        12'h0AC: sinewave <= 12'h215;
        12'h0AD: sinewave <= 12'h218;
        12'h0AE: sinewave <= 12'h21B;
        12'h0AF: sinewave <= 12'h21E;
        12'h0B0: sinewave <= 12'h221;
        12'h0B1: sinewave <= 12'h224;
        12'h0B2: sinewave <= 12'h228;
        12'h0B3: sinewave <= 12'h22B;
        12'h0B4: sinewave <= 12'h22E;
        12'h0B5: sinewave <= 12'h231;
        12'h0B6: sinewave <= 12'h234;
        12'h0B7: sinewave <= 12'h237;
        12'h0B8: sinewave <= 12'h23A;
        12'h0B9: sinewave <= 12'h23D;
        12'h0BA: sinewave <= 12'h240;
        12'h0BB: sinewave <= 12'h243;
        12'h0BC: sinewave <= 12'h246;
        12'h0BD: sinewave <= 12'h249;
        12'h0BE: sinewave <= 12'h24C;
        12'h0BF: sinewave <= 12'h24F;
        12'h0C0: sinewave <= 12'h252;
        12'h0C1: sinewave <= 12'h255;
        12'h0C2: sinewave <= 12'h258;
        12'h0C3: sinewave <= 12'h25B;
        12'h0C4: sinewave <= 12'h25E;
        12'h0C5: sinewave <= 12'h261;
        12'h0C6: sinewave <= 12'h264;
        12'h0C7: sinewave <= 12'h267;
        12'h0C8: sinewave <= 12'h26A;
        12'h0C9: sinewave <= 12'h26D;
        12'h0CA: sinewave <= 12'h270;
        12'h0CB: sinewave <= 12'h273;
        12'h0CC: sinewave <= 12'h276;
        12'h0CD: sinewave <= 12'h279;
        12'h0CE: sinewave <= 12'h27C;
        12'h0CF: sinewave <= 12'h27F;
        12'h0D0: sinewave <= 12'h282;
        12'h0D1: sinewave <= 12'h285;
        12'h0D2: sinewave <= 12'h288;
        12'h0D3: sinewave <= 12'h28B;
        12'h0D4: sinewave <= 12'h28E;
        12'h0D5: sinewave <= 12'h290;
        12'h0D6: sinewave <= 12'h293;
        12'h0D7: sinewave <= 12'h296;
        12'h0D8: sinewave <= 12'h299;
        12'h0D9: sinewave <= 12'h29C;
        12'h0DA: sinewave <= 12'h29F;
        12'h0DB: sinewave <= 12'h2A2;
        12'h0DC: sinewave <= 12'h2A5;
        12'h0DD: sinewave <= 12'h2A8;
        12'h0DE: sinewave <= 12'h2AB;
        12'h0DF: sinewave <= 12'h2AE;
        12'h0E0: sinewave <= 12'h2B1;
        12'h0E1: sinewave <= 12'h2B4;
        12'h0E2: sinewave <= 12'h2B7;
        12'h0E3: sinewave <= 12'h2BA;
        12'h0E4: sinewave <= 12'h2BD;
        12'h0E5: sinewave <= 12'h2C0;
        12'h0E6: sinewave <= 12'h2C3;
        12'h0E7: sinewave <= 12'h2C6;
        12'h0E8: sinewave <= 12'h2C9;
        12'h0E9: sinewave <= 12'h2CC;
        12'h0EA: sinewave <= 12'h2CF;
        12'h0EB: sinewave <= 12'h2D2;
        12'h0EC: sinewave <= 12'h2D4;
        12'h0ED: sinewave <= 12'h2D7;
        12'h0EE: sinewave <= 12'h2DA;
        12'h0EF: sinewave <= 12'h2DD;
        12'h0F0: sinewave <= 12'h2E0;
        12'h0F1: sinewave <= 12'h2E3;
        12'h0F2: sinewave <= 12'h2E6;
        12'h0F3: sinewave <= 12'h2E9;
        12'h0F4: sinewave <= 12'h2EC;
        12'h0F5: sinewave <= 12'h2EF;
        12'h0F6: sinewave <= 12'h2F2;
        12'h0F7: sinewave <= 12'h2F5;
        12'h0F8: sinewave <= 12'h2F8;
        12'h0F9: sinewave <= 12'h2FB;
        12'h0FA: sinewave <= 12'h2FD;
        12'h0FB: sinewave <= 12'h300;
        12'h0FC: sinewave <= 12'h303;
        12'h0FD: sinewave <= 12'h306;
        12'h0FE: sinewave <= 12'h309;
        12'h0FF: sinewave <= 12'h30C;
        12'h100: sinewave <= 12'h30F;
        12'h101: sinewave <= 12'h312;
        12'h102: sinewave <= 12'h315;
        12'h103: sinewave <= 12'h318;
        12'h104: sinewave <= 12'h31A;
        12'h105: sinewave <= 12'h31D;
        12'h106: sinewave <= 12'h320;
        12'h107: sinewave <= 12'h323;
        12'h108: sinewave <= 12'h326;
        12'h109: sinewave <= 12'h329;
        12'h10A: sinewave <= 12'h32C;
        12'h10B: sinewave <= 12'h32F;
        12'h10C: sinewave <= 12'h332;
        12'h10D: sinewave <= 12'h334;
        12'h10E: sinewave <= 12'h337;
        12'h10F: sinewave <= 12'h33A;
        12'h110: sinewave <= 12'h33D;
        12'h111: sinewave <= 12'h340;
        12'h112: sinewave <= 12'h343;
        12'h113: sinewave <= 12'h346;
        12'h114: sinewave <= 12'h348;
        12'h115: sinewave <= 12'h34B;
        12'h116: sinewave <= 12'h34E;
        12'h117: sinewave <= 12'h351;
        12'h118: sinewave <= 12'h354;
        12'h119: sinewave <= 12'h357;
        12'h11A: sinewave <= 12'h35A;
        12'h11B: sinewave <= 12'h35C;
        12'h11C: sinewave <= 12'h35F;
        12'h11D: sinewave <= 12'h362;
        12'h11E: sinewave <= 12'h365;
        12'h11F: sinewave <= 12'h368;
        12'h120: sinewave <= 12'h36B;
        12'h121: sinewave <= 12'h36E;
        12'h122: sinewave <= 12'h370;
        12'h123: sinewave <= 12'h373;
        12'h124: sinewave <= 12'h376;
        12'h125: sinewave <= 12'h379;
        12'h126: sinewave <= 12'h37C;
        12'h127: sinewave <= 12'h37F;
        12'h128: sinewave <= 12'h381;
        12'h129: sinewave <= 12'h384;
        12'h12A: sinewave <= 12'h387;
        12'h12B: sinewave <= 12'h38A;
        12'h12C: sinewave <= 12'h38D;
        12'h12D: sinewave <= 12'h38F;
        12'h12E: sinewave <= 12'h392;
        12'h12F: sinewave <= 12'h395;
        12'h130: sinewave <= 12'h398;
        12'h131: sinewave <= 12'h39B;
        12'h132: sinewave <= 12'h39D;
        12'h133: sinewave <= 12'h3A0;
        12'h134: sinewave <= 12'h3A3;
        12'h135: sinewave <= 12'h3A6;
        12'h136: sinewave <= 12'h3A9;
        12'h137: sinewave <= 12'h3AB;
        12'h138: sinewave <= 12'h3AE;
        12'h139: sinewave <= 12'h3B1;
        12'h13A: sinewave <= 12'h3B4;
        12'h13B: sinewave <= 12'h3B7;
        12'h13C: sinewave <= 12'h3B9;
        12'h13D: sinewave <= 12'h3BC;
        12'h13E: sinewave <= 12'h3BF;
        12'h13F: sinewave <= 12'h3C2;
        12'h140: sinewave <= 12'h3C4;
        12'h141: sinewave <= 12'h3C7;
        12'h142: sinewave <= 12'h3CA;
        12'h143: sinewave <= 12'h3CD;
        12'h144: sinewave <= 12'h3D0;
        12'h145: sinewave <= 12'h3D2;
        12'h146: sinewave <= 12'h3D5;
        12'h147: sinewave <= 12'h3D8;
        12'h148: sinewave <= 12'h3DB;
        12'h149: sinewave <= 12'h3DD;
        12'h14A: sinewave <= 12'h3E0;
        12'h14B: sinewave <= 12'h3E3;
        12'h14C: sinewave <= 12'h3E6;
        12'h14D: sinewave <= 12'h3E8;
        12'h14E: sinewave <= 12'h3EB;
        12'h14F: sinewave <= 12'h3EE;
        12'h150: sinewave <= 12'h3F0;
        12'h151: sinewave <= 12'h3F3;
        12'h152: sinewave <= 12'h3F6;
        12'h153: sinewave <= 12'h3F9;
        12'h154: sinewave <= 12'h3FB;
        12'h155: sinewave <= 12'h3FE;
        12'h156: sinewave <= 12'h401;
        12'h157: sinewave <= 12'h404;
        12'h158: sinewave <= 12'h406;
        12'h159: sinewave <= 12'h409;
        12'h15A: sinewave <= 12'h40C;
        12'h15B: sinewave <= 12'h40E;
        12'h15C: sinewave <= 12'h411;
        12'h15D: sinewave <= 12'h414;
        12'h15E: sinewave <= 12'h416;
        12'h15F: sinewave <= 12'h419;
        12'h160: sinewave <= 12'h41C;
        12'h161: sinewave <= 12'h41F;
        12'h162: sinewave <= 12'h421;
        12'h163: sinewave <= 12'h424;
        12'h164: sinewave <= 12'h427;
        12'h165: sinewave <= 12'h429;
        12'h166: sinewave <= 12'h42C;
        12'h167: sinewave <= 12'h42F;
        12'h168: sinewave <= 12'h431;
        12'h169: sinewave <= 12'h434;
        12'h16A: sinewave <= 12'h437;
        12'h16B: sinewave <= 12'h439;
        12'h16C: sinewave <= 12'h43C;
        12'h16D: sinewave <= 12'h43F;
        12'h16E: sinewave <= 12'h441;
        12'h16F: sinewave <= 12'h444;
        12'h170: sinewave <= 12'h447;
        12'h171: sinewave <= 12'h449;
        12'h172: sinewave <= 12'h44C;
        12'h173: sinewave <= 12'h44F;
        12'h174: sinewave <= 12'h451;
        12'h175: sinewave <= 12'h454;
        12'h176: sinewave <= 12'h457;
        12'h177: sinewave <= 12'h459;
        12'h178: sinewave <= 12'h45C;
        12'h179: sinewave <= 12'h45E;
        12'h17A: sinewave <= 12'h461;
        12'h17B: sinewave <= 12'h464;
        12'h17C: sinewave <= 12'h466;
        12'h17D: sinewave <= 12'h469;
        12'h17E: sinewave <= 12'h46C;
        12'h17F: sinewave <= 12'h46E;
        12'h180: sinewave <= 12'h471;
        12'h181: sinewave <= 12'h473;
        12'h182: sinewave <= 12'h476;
        12'h183: sinewave <= 12'h479;
        12'h184: sinewave <= 12'h47B;
        12'h185: sinewave <= 12'h47E;
        12'h186: sinewave <= 12'h480;
        12'h187: sinewave <= 12'h483;
        12'h188: sinewave <= 12'h486;
        12'h189: sinewave <= 12'h488;
        12'h18A: sinewave <= 12'h48B;
        12'h18B: sinewave <= 12'h48D;
        12'h18C: sinewave <= 12'h490;
        12'h18D: sinewave <= 12'h492;
        12'h18E: sinewave <= 12'h495;
        12'h18F: sinewave <= 12'h498;
        12'h190: sinewave <= 12'h49A;
        12'h191: sinewave <= 12'h49D;
        12'h192: sinewave <= 12'h49F;
        12'h193: sinewave <= 12'h4A2;
        12'h194: sinewave <= 12'h4A4;
        12'h195: sinewave <= 12'h4A7;
        12'h196: sinewave <= 12'h4AA;
        12'h197: sinewave <= 12'h4AC;
        12'h198: sinewave <= 12'h4AF;
        12'h199: sinewave <= 12'h4B1;
        12'h19A: sinewave <= 12'h4B4;
        12'h19B: sinewave <= 12'h4B6;
        12'h19C: sinewave <= 12'h4B9;
        12'h19D: sinewave <= 12'h4BB;
        12'h19E: sinewave <= 12'h4BE;
        12'h19F: sinewave <= 12'h4C0;
        12'h1A0: sinewave <= 12'h4C3;
        12'h1A1: sinewave <= 12'h4C5;
        12'h1A2: sinewave <= 12'h4C8;
        12'h1A3: sinewave <= 12'h4CA;
        12'h1A4: sinewave <= 12'h4CD;
        12'h1A5: sinewave <= 12'h4CF;
        12'h1A6: sinewave <= 12'h4D2;
        12'h1A7: sinewave <= 12'h4D4;
        12'h1A8: sinewave <= 12'h4D7;
        12'h1A9: sinewave <= 12'h4D9;
        12'h1AA: sinewave <= 12'h4DC;
        12'h1AB: sinewave <= 12'h4DE;
        12'h1AC: sinewave <= 12'h4E1;
        12'h1AD: sinewave <= 12'h4E3;
        12'h1AE: sinewave <= 12'h4E6;
        12'h1AF: sinewave <= 12'h4E8;
        12'h1B0: sinewave <= 12'h4EB;
        12'h1B1: sinewave <= 12'h4ED;
        12'h1B2: sinewave <= 12'h4F0;
        12'h1B3: sinewave <= 12'h4F2;
        12'h1B4: sinewave <= 12'h4F5;
        12'h1B5: sinewave <= 12'h4F7;
        12'h1B6: sinewave <= 12'h4FA;
        12'h1B7: sinewave <= 12'h4FC;
        12'h1B8: sinewave <= 12'h4FF;
        12'h1B9: sinewave <= 12'h501;
        12'h1BA: sinewave <= 12'h503;
        12'h1BB: sinewave <= 12'h506;
        12'h1BC: sinewave <= 12'h508;
        12'h1BD: sinewave <= 12'h50B;
        12'h1BE: sinewave <= 12'h50D;
        12'h1BF: sinewave <= 12'h510;
        12'h1C0: sinewave <= 12'h512;
        12'h1C1: sinewave <= 12'h515;
        12'h1C2: sinewave <= 12'h517;
        12'h1C3: sinewave <= 12'h519;
        12'h1C4: sinewave <= 12'h51C;
        12'h1C5: sinewave <= 12'h51E;
        12'h1C6: sinewave <= 12'h521;
        12'h1C7: sinewave <= 12'h523;
        12'h1C8: sinewave <= 12'h525;
        12'h1C9: sinewave <= 12'h528;
        12'h1CA: sinewave <= 12'h52A;
        12'h1CB: sinewave <= 12'h52D;
        12'h1CC: sinewave <= 12'h52F;
        12'h1CD: sinewave <= 12'h531;
        12'h1CE: sinewave <= 12'h534;
        12'h1CF: sinewave <= 12'h536;
        12'h1D0: sinewave <= 12'h539;
        12'h1D1: sinewave <= 12'h53B;
        12'h1D2: sinewave <= 12'h53D;
        12'h1D3: sinewave <= 12'h540;
        12'h1D4: sinewave <= 12'h542;
        12'h1D5: sinewave <= 12'h544;
        12'h1D6: sinewave <= 12'h547;
        12'h1D7: sinewave <= 12'h549;
        12'h1D8: sinewave <= 12'h54B;
        12'h1D9: sinewave <= 12'h54E;
        12'h1DA: sinewave <= 12'h550;
        12'h1DB: sinewave <= 12'h553;
        12'h1DC: sinewave <= 12'h555;
        12'h1DD: sinewave <= 12'h557;
        12'h1DE: sinewave <= 12'h55A;
        12'h1DF: sinewave <= 12'h55C;
        12'h1E0: sinewave <= 12'h55E;
        12'h1E1: sinewave <= 12'h561;
        12'h1E2: sinewave <= 12'h563;
        12'h1E3: sinewave <= 12'h565;
        12'h1E4: sinewave <= 12'h567;
        12'h1E5: sinewave <= 12'h56A;
        12'h1E6: sinewave <= 12'h56C;
        12'h1E7: sinewave <= 12'h56E;
        12'h1E8: sinewave <= 12'h571;
        12'h1E9: sinewave <= 12'h573;
        12'h1EA: sinewave <= 12'h575;
        12'h1EB: sinewave <= 12'h578;
        12'h1EC: sinewave <= 12'h57A;
        12'h1ED: sinewave <= 12'h57C;
        12'h1EE: sinewave <= 12'h57E;
        12'h1EF: sinewave <= 12'h581;
        12'h1F0: sinewave <= 12'h583;
        12'h1F1: sinewave <= 12'h585;
        12'h1F2: sinewave <= 12'h588;
        12'h1F3: sinewave <= 12'h58A;
        12'h1F4: sinewave <= 12'h58C;
        12'h1F5: sinewave <= 12'h58E;
        12'h1F6: sinewave <= 12'h591;
        12'h1F7: sinewave <= 12'h593;
        12'h1F8: sinewave <= 12'h595;
        12'h1F9: sinewave <= 12'h597;
        12'h1FA: sinewave <= 12'h59A;
        12'h1FB: sinewave <= 12'h59C;
        12'h1FC: sinewave <= 12'h59E;
        12'h1FD: sinewave <= 12'h5A0;
        12'h1FE: sinewave <= 12'h5A3;
        12'h1FF: sinewave <= 12'h5A5;
        12'h200: sinewave <= 12'h5A7;
        12'h201: sinewave <= 12'h5A9;
        12'h202: sinewave <= 12'h5AB;
        12'h203: sinewave <= 12'h5AE;
        12'h204: sinewave <= 12'h5B0;
        12'h205: sinewave <= 12'h5B2;
        12'h206: sinewave <= 12'h5B4;
        12'h207: sinewave <= 12'h5B6;
        12'h208: sinewave <= 12'h5B9;
        12'h209: sinewave <= 12'h5BB;
        12'h20A: sinewave <= 12'h5BD;
        12'h20B: sinewave <= 12'h5BF;
        12'h20C: sinewave <= 12'h5C1;
        12'h20D: sinewave <= 12'h5C4;
        12'h20E: sinewave <= 12'h5C6;
        12'h20F: sinewave <= 12'h5C8;
        12'h210: sinewave <= 12'h5CA;
        12'h211: sinewave <= 12'h5CC;
        12'h212: sinewave <= 12'h5CE;
        12'h213: sinewave <= 12'h5D1;
        12'h214: sinewave <= 12'h5D3;
        12'h215: sinewave <= 12'h5D5;
        12'h216: sinewave <= 12'h5D7;
        12'h217: sinewave <= 12'h5D9;
        12'h218: sinewave <= 12'h5DB;
        12'h219: sinewave <= 12'h5DD;
        12'h21A: sinewave <= 12'h5E0;
        12'h21B: sinewave <= 12'h5E2;
        12'h21C: sinewave <= 12'h5E4;
        12'h21D: sinewave <= 12'h5E6;
        12'h21E: sinewave <= 12'h5E8;
        12'h21F: sinewave <= 12'h5EA;
        12'h220: sinewave <= 12'h5EC;
        12'h221: sinewave <= 12'h5EE;
        12'h222: sinewave <= 12'h5F0;
        12'h223: sinewave <= 12'h5F3;
        12'h224: sinewave <= 12'h5F5;
        12'h225: sinewave <= 12'h5F7;
        12'h226: sinewave <= 12'h5F9;
        12'h227: sinewave <= 12'h5FB;
        12'h228: sinewave <= 12'h5FD;
        12'h229: sinewave <= 12'h5FF;
        12'h22A: sinewave <= 12'h601;
        12'h22B: sinewave <= 12'h603;
        12'h22C: sinewave <= 12'h605;
        12'h22D: sinewave <= 12'h607;
        12'h22E: sinewave <= 12'h609;
        12'h22F: sinewave <= 12'h60B;
        12'h230: sinewave <= 12'h60E;
        12'h231: sinewave <= 12'h610;
        12'h232: sinewave <= 12'h612;
        12'h233: sinewave <= 12'h614;
        12'h234: sinewave <= 12'h616;
        12'h235: sinewave <= 12'h618;
        12'h236: sinewave <= 12'h61A;
        12'h237: sinewave <= 12'h61C;
        12'h238: sinewave <= 12'h61E;
        12'h239: sinewave <= 12'h620;
        12'h23A: sinewave <= 12'h622;
        12'h23B: sinewave <= 12'h624;
        12'h23C: sinewave <= 12'h626;
        12'h23D: sinewave <= 12'h628;
        12'h23E: sinewave <= 12'h62A;
        12'h23F: sinewave <= 12'h62C;
        12'h240: sinewave <= 12'h62E;
        12'h241: sinewave <= 12'h630;
        12'h242: sinewave <= 12'h632;
        12'h243: sinewave <= 12'h634;
        12'h244: sinewave <= 12'h636;
        12'h245: sinewave <= 12'h638;
        12'h246: sinewave <= 12'h63A;
        12'h247: sinewave <= 12'h63C;
        12'h248: sinewave <= 12'h63E;
        12'h249: sinewave <= 12'h640;
        12'h24A: sinewave <= 12'h642;
        12'h24B: sinewave <= 12'h644;
        12'h24C: sinewave <= 12'h645;
        12'h24D: sinewave <= 12'h647;
        12'h24E: sinewave <= 12'h649;
        12'h24F: sinewave <= 12'h64B;
        12'h250: sinewave <= 12'h64D;
        12'h251: sinewave <= 12'h64F;
        12'h252: sinewave <= 12'h651;
        12'h253: sinewave <= 12'h653;
        12'h254: sinewave <= 12'h655;
        12'h255: sinewave <= 12'h657;
        12'h256: sinewave <= 12'h659;
        12'h257: sinewave <= 12'h65B;
        12'h258: sinewave <= 12'h65D;
        12'h259: sinewave <= 12'h65E;
        12'h25A: sinewave <= 12'h660;
        12'h25B: sinewave <= 12'h662;
        12'h25C: sinewave <= 12'h664;
        12'h25D: sinewave <= 12'h666;
        12'h25E: sinewave <= 12'h668;
        12'h25F: sinewave <= 12'h66A;
        12'h260: sinewave <= 12'h66C;
        12'h261: sinewave <= 12'h66E;
        12'h262: sinewave <= 12'h66F;
        12'h263: sinewave <= 12'h671;
        12'h264: sinewave <= 12'h673;
        12'h265: sinewave <= 12'h675;
        12'h266: sinewave <= 12'h677;
        12'h267: sinewave <= 12'h679;
        12'h268: sinewave <= 12'h67B;
        12'h269: sinewave <= 12'h67C;
        12'h26A: sinewave <= 12'h67E;
        12'h26B: sinewave <= 12'h680;
        12'h26C: sinewave <= 12'h682;
        12'h26D: sinewave <= 12'h684;
        12'h26E: sinewave <= 12'h685;
        12'h26F: sinewave <= 12'h687;
        12'h270: sinewave <= 12'h689;
        12'h271: sinewave <= 12'h68B;
        12'h272: sinewave <= 12'h68D;
        12'h273: sinewave <= 12'h68F;
        12'h274: sinewave <= 12'h690;
        12'h275: sinewave <= 12'h692;
        12'h276: sinewave <= 12'h694;
        12'h277: sinewave <= 12'h696;
        12'h278: sinewave <= 12'h697;
        12'h279: sinewave <= 12'h699;
        12'h27A: sinewave <= 12'h69B;
        12'h27B: sinewave <= 12'h69D;
        12'h27C: sinewave <= 12'h69F;
        12'h27D: sinewave <= 12'h6A0;
        12'h27E: sinewave <= 12'h6A2;
        12'h27F: sinewave <= 12'h6A4;
        12'h280: sinewave <= 12'h6A6;
        12'h281: sinewave <= 12'h6A7;
        12'h282: sinewave <= 12'h6A9;
        12'h283: sinewave <= 12'h6AB;
        12'h284: sinewave <= 12'h6AC;
        12'h285: sinewave <= 12'h6AE;
        12'h286: sinewave <= 12'h6B0;
        12'h287: sinewave <= 12'h6B2;
        12'h288: sinewave <= 12'h6B3;
        12'h289: sinewave <= 12'h6B5;
        12'h28A: sinewave <= 12'h6B7;
        12'h28B: sinewave <= 12'h6B8;
        12'h28C: sinewave <= 12'h6BA;
        12'h28D: sinewave <= 12'h6BC;
        12'h28E: sinewave <= 12'h6BE;
        12'h28F: sinewave <= 12'h6BF;
        12'h290: sinewave <= 12'h6C1;
        12'h291: sinewave <= 12'h6C3;
        12'h292: sinewave <= 12'h6C4;
        12'h293: sinewave <= 12'h6C6;
        12'h294: sinewave <= 12'h6C8;
        12'h295: sinewave <= 12'h6C9;
        12'h296: sinewave <= 12'h6CB;
        12'h297: sinewave <= 12'h6CD;
        12'h298: sinewave <= 12'h6CE;
        12'h299: sinewave <= 12'h6D0;
        12'h29A: sinewave <= 12'h6D2;
        12'h29B: sinewave <= 12'h6D3;
        12'h29C: sinewave <= 12'h6D5;
        12'h29D: sinewave <= 12'h6D6;
        12'h29E: sinewave <= 12'h6D8;
        12'h29F: sinewave <= 12'h6DA;
        12'h2A0: sinewave <= 12'h6DB;
        12'h2A1: sinewave <= 12'h6DD;
        12'h2A2: sinewave <= 12'h6DE;
        12'h2A3: sinewave <= 12'h6E0;
        12'h2A4: sinewave <= 12'h6E2;
        12'h2A5: sinewave <= 12'h6E3;
        12'h2A6: sinewave <= 12'h6E5;
        12'h2A7: sinewave <= 12'h6E6;
        12'h2A8: sinewave <= 12'h6E8;
        12'h2A9: sinewave <= 12'h6EA;
        12'h2AA: sinewave <= 12'h6EB;
        12'h2AB: sinewave <= 12'h6ED;
        12'h2AC: sinewave <= 12'h6EE;
        12'h2AD: sinewave <= 12'h6F0;
        12'h2AE: sinewave <= 12'h6F1;
        12'h2AF: sinewave <= 12'h6F3;
        12'h2B0: sinewave <= 12'h6F5;
        12'h2B1: sinewave <= 12'h6F6;
        12'h2B2: sinewave <= 12'h6F8;
        12'h2B3: sinewave <= 12'h6F9;
        12'h2B4: sinewave <= 12'h6FB;
        12'h2B5: sinewave <= 12'h6FC;
        12'h2B6: sinewave <= 12'h6FE;
        12'h2B7: sinewave <= 12'h6FF;
        12'h2B8: sinewave <= 12'h701;
        12'h2B9: sinewave <= 12'h702;
        12'h2BA: sinewave <= 12'h704;
        12'h2BB: sinewave <= 12'h705;
        12'h2BC: sinewave <= 12'h707;
        12'h2BD: sinewave <= 12'h708;
        12'h2BE: sinewave <= 12'h70A;
        12'h2BF: sinewave <= 12'h70B;
        12'h2C0: sinewave <= 12'h70D;
        12'h2C1: sinewave <= 12'h70E;
        12'h2C2: sinewave <= 12'h710;
        12'h2C3: sinewave <= 12'h711;
        12'h2C4: sinewave <= 12'h713;
        12'h2C5: sinewave <= 12'h714;
        12'h2C6: sinewave <= 12'h716;
        12'h2C7: sinewave <= 12'h717;
        12'h2C8: sinewave <= 12'h718;
        12'h2C9: sinewave <= 12'h71A;
        12'h2CA: sinewave <= 12'h71B;
        12'h2CB: sinewave <= 12'h71D;
        12'h2CC: sinewave <= 12'h71E;
        12'h2CD: sinewave <= 12'h720;
        12'h2CE: sinewave <= 12'h721;
        12'h2CF: sinewave <= 12'h723;
        12'h2D0: sinewave <= 12'h724;
        12'h2D1: sinewave <= 12'h725;
        12'h2D2: sinewave <= 12'h727;
        12'h2D3: sinewave <= 12'h728;
        12'h2D4: sinewave <= 12'h72A;
        12'h2D5: sinewave <= 12'h72B;
        12'h2D6: sinewave <= 12'h72C;
        12'h2D7: sinewave <= 12'h72E;
        12'h2D8: sinewave <= 12'h72F;
        12'h2D9: sinewave <= 12'h730;
        12'h2DA: sinewave <= 12'h732;
        12'h2DB: sinewave <= 12'h733;
        12'h2DC: sinewave <= 12'h735;
        12'h2DD: sinewave <= 12'h736;
        12'h2DE: sinewave <= 12'h737;
        12'h2DF: sinewave <= 12'h739;
        12'h2E0: sinewave <= 12'h73A;
        12'h2E1: sinewave <= 12'h73B;
        12'h2E2: sinewave <= 12'h73D;
        12'h2E3: sinewave <= 12'h73E;
        12'h2E4: sinewave <= 12'h73F;
        12'h2E5: sinewave <= 12'h741;
        12'h2E6: sinewave <= 12'h742;
        12'h2E7: sinewave <= 12'h743;
        12'h2E8: sinewave <= 12'h745;
        12'h2E9: sinewave <= 12'h746;
        12'h2EA: sinewave <= 12'h747;
        12'h2EB: sinewave <= 12'h748;
        12'h2EC: sinewave <= 12'h74A;
        12'h2ED: sinewave <= 12'h74B;
        12'h2EE: sinewave <= 12'h74C;
        12'h2EF: sinewave <= 12'h74E;
        12'h2F0: sinewave <= 12'h74F;
        12'h2F1: sinewave <= 12'h750;
        12'h2F2: sinewave <= 12'h751;
        12'h2F3: sinewave <= 12'h753;
        12'h2F4: sinewave <= 12'h754;
        12'h2F5: sinewave <= 12'h755;
        12'h2F6: sinewave <= 12'h756;
        12'h2F7: sinewave <= 12'h758;
        12'h2F8: sinewave <= 12'h759;
        12'h2F9: sinewave <= 12'h75A;
        12'h2FA: sinewave <= 12'h75B;
        12'h2FB: sinewave <= 12'h75D;
        12'h2FC: sinewave <= 12'h75E;
        12'h2FD: sinewave <= 12'h75F;
        12'h2FE: sinewave <= 12'h760;
        12'h2FF: sinewave <= 12'h761;
        12'h300: sinewave <= 12'h763;
        12'h301: sinewave <= 12'h764;
        12'h302: sinewave <= 12'h765;
        12'h303: sinewave <= 12'h766;
        12'h304: sinewave <= 12'h767;
        12'h305: sinewave <= 12'h769;
        12'h306: sinewave <= 12'h76A;
        12'h307: sinewave <= 12'h76B;
        12'h308: sinewave <= 12'h76C;
        12'h309: sinewave <= 12'h76D;
        12'h30A: sinewave <= 12'h76E;
        12'h30B: sinewave <= 12'h770;
        12'h30C: sinewave <= 12'h771;
        12'h30D: sinewave <= 12'h772;
        12'h30E: sinewave <= 12'h773;
        12'h30F: sinewave <= 12'h774;
        12'h310: sinewave <= 12'h775;
        12'h311: sinewave <= 12'h776;
        12'h312: sinewave <= 12'h778;
        12'h313: sinewave <= 12'h779;
        12'h314: sinewave <= 12'h77A;
        12'h315: sinewave <= 12'h77B;
        12'h316: sinewave <= 12'h77C;
        12'h317: sinewave <= 12'h77D;
        12'h318: sinewave <= 12'h77E;
        12'h319: sinewave <= 12'h77F;
        12'h31A: sinewave <= 12'h780;
        12'h31B: sinewave <= 12'h781;
        12'h31C: sinewave <= 12'h783;
        12'h31D: sinewave <= 12'h784;
        12'h31E: sinewave <= 12'h785;
        12'h31F: sinewave <= 12'h786;
        12'h320: sinewave <= 12'h787;
        12'h321: sinewave <= 12'h788;
        12'h322: sinewave <= 12'h789;
        12'h323: sinewave <= 12'h78A;
        12'h324: sinewave <= 12'h78B;
        12'h325: sinewave <= 12'h78C;
        12'h326: sinewave <= 12'h78D;
        12'h327: sinewave <= 12'h78E;
        12'h328: sinewave <= 12'h78F;
        12'h329: sinewave <= 12'h790;
        12'h32A: sinewave <= 12'h791;
        12'h32B: sinewave <= 12'h792;
        12'h32C: sinewave <= 12'h793;
        12'h32D: sinewave <= 12'h794;
        12'h32E: sinewave <= 12'h795;
        12'h32F: sinewave <= 12'h796;
        12'h330: sinewave <= 12'h797;
        12'h331: sinewave <= 12'h798;
        12'h332: sinewave <= 12'h799;
        12'h333: sinewave <= 12'h79A;
        12'h334: sinewave <= 12'h79B;
        12'h335: sinewave <= 12'h79C;
        12'h336: sinewave <= 12'h79D;
        12'h337: sinewave <= 12'h79E;
        12'h338: sinewave <= 12'h79F;
        12'h339: sinewave <= 12'h7A0;
        12'h33A: sinewave <= 12'h7A1;
        12'h33B: sinewave <= 12'h7A2;
        12'h33C: sinewave <= 12'h7A3;
        12'h33D: sinewave <= 12'h7A4;
        12'h33E: sinewave <= 12'h7A5;
        12'h33F: sinewave <= 12'h7A5;
        12'h340: sinewave <= 12'h7A6;
        12'h341: sinewave <= 12'h7A7;
        12'h342: sinewave <= 12'h7A8;
        12'h343: sinewave <= 12'h7A9;
        12'h344: sinewave <= 12'h7AA;
        12'h345: sinewave <= 12'h7AB;
        12'h346: sinewave <= 12'h7AC;
        12'h347: sinewave <= 12'h7AD;
        12'h348: sinewave <= 12'h7AE;
        12'h349: sinewave <= 12'h7AE;
        12'h34A: sinewave <= 12'h7AF;
        12'h34B: sinewave <= 12'h7B0;
        12'h34C: sinewave <= 12'h7B1;
        12'h34D: sinewave <= 12'h7B2;
        12'h34E: sinewave <= 12'h7B3;
        12'h34F: sinewave <= 12'h7B4;
        12'h350: sinewave <= 12'h7B4;
        12'h351: sinewave <= 12'h7B5;
        12'h352: sinewave <= 12'h7B6;
        12'h353: sinewave <= 12'h7B7;
        12'h354: sinewave <= 12'h7B8;
        12'h355: sinewave <= 12'h7B8;
        12'h356: sinewave <= 12'h7B9;
        12'h357: sinewave <= 12'h7BA;
        12'h358: sinewave <= 12'h7BB;
        12'h359: sinewave <= 12'h7BC;
        12'h35A: sinewave <= 12'h7BC;
        12'h35B: sinewave <= 12'h7BD;
        12'h35C: sinewave <= 12'h7BE;
        12'h35D: sinewave <= 12'h7BF;
        12'h35E: sinewave <= 12'h7C0;
        12'h35F: sinewave <= 12'h7C0;
        12'h360: sinewave <= 12'h7C1;
        12'h361: sinewave <= 12'h7C2;
        12'h362: sinewave <= 12'h7C3;
        12'h363: sinewave <= 12'h7C3;
        12'h364: sinewave <= 12'h7C4;
        12'h365: sinewave <= 12'h7C5;
        12'h366: sinewave <= 12'h7C6;
        12'h367: sinewave <= 12'h7C6;
        12'h368: sinewave <= 12'h7C7;
        12'h369: sinewave <= 12'h7C8;
        12'h36A: sinewave <= 12'h7C9;
        12'h36B: sinewave <= 12'h7C9;
        12'h36C: sinewave <= 12'h7CA;
        12'h36D: sinewave <= 12'h7CB;
        12'h36E: sinewave <= 12'h7CB;
        12'h36F: sinewave <= 12'h7CC;
        12'h370: sinewave <= 12'h7CD;
        12'h371: sinewave <= 12'h7CD;
        12'h372: sinewave <= 12'h7CE;
        12'h373: sinewave <= 12'h7CF;
        12'h374: sinewave <= 12'h7CF;
        12'h375: sinewave <= 12'h7D0;
        12'h376: sinewave <= 12'h7D1;
        12'h377: sinewave <= 12'h7D1;
        12'h378: sinewave <= 12'h7D2;
        12'h379: sinewave <= 12'h7D3;
        12'h37A: sinewave <= 12'h7D3;
        12'h37B: sinewave <= 12'h7D4;
        12'h37C: sinewave <= 12'h7D5;
        12'h37D: sinewave <= 12'h7D5;
        12'h37E: sinewave <= 12'h7D6;
        12'h37F: sinewave <= 12'h7D7;
        12'h380: sinewave <= 12'h7D7;
        12'h381: sinewave <= 12'h7D8;
        12'h382: sinewave <= 12'h7D8;
        12'h383: sinewave <= 12'h7D9;
        12'h384: sinewave <= 12'h7DA;
        12'h385: sinewave <= 12'h7DA;
        12'h386: sinewave <= 12'h7DB;
        12'h387: sinewave <= 12'h7DB;
        12'h388: sinewave <= 12'h7DC;
        12'h389: sinewave <= 12'h7DC;
        12'h38A: sinewave <= 12'h7DD;
        12'h38B: sinewave <= 12'h7DE;
        12'h38C: sinewave <= 12'h7DE;
        12'h38D: sinewave <= 12'h7DF;
        12'h38E: sinewave <= 12'h7DF;
        12'h38F: sinewave <= 12'h7E0;
        12'h390: sinewave <= 12'h7E0;
        12'h391: sinewave <= 12'h7E1;
        12'h392: sinewave <= 12'h7E1;
        12'h393: sinewave <= 12'h7E2;
        12'h394: sinewave <= 12'h7E2;
        12'h395: sinewave <= 12'h7E3;
        12'h396: sinewave <= 12'h7E3;
        12'h397: sinewave <= 12'h7E4;
        12'h398: sinewave <= 12'h7E5;
        12'h399: sinewave <= 12'h7E5;
        12'h39A: sinewave <= 12'h7E5;
        12'h39B: sinewave <= 12'h7E6;
        12'h39C: sinewave <= 12'h7E6;
        12'h39D: sinewave <= 12'h7E7;
        12'h39E: sinewave <= 12'h7E7;
        12'h39F: sinewave <= 12'h7E8;
        12'h3A0: sinewave <= 12'h7E8;
        12'h3A1: sinewave <= 12'h7E9;
        12'h3A2: sinewave <= 12'h7E9;
        12'h3A3: sinewave <= 12'h7EA;
        12'h3A4: sinewave <= 12'h7EA;
        12'h3A5: sinewave <= 12'h7EB;
        12'h3A6: sinewave <= 12'h7EB;
        12'h3A7: sinewave <= 12'h7EB;
        12'h3A8: sinewave <= 12'h7EC;
        12'h3A9: sinewave <= 12'h7EC;
        12'h3AA: sinewave <= 12'h7ED;
        12'h3AB: sinewave <= 12'h7ED;
        12'h3AC: sinewave <= 12'h7EE;
        12'h3AD: sinewave <= 12'h7EE;
        12'h3AE: sinewave <= 12'h7EE;
        12'h3AF: sinewave <= 12'h7EF;
        12'h3B0: sinewave <= 12'h7EF;
        12'h3B1: sinewave <= 12'h7EF;
        12'h3B2: sinewave <= 12'h7F0;
        12'h3B3: sinewave <= 12'h7F0;
        12'h3B4: sinewave <= 12'h7F1;
        12'h3B5: sinewave <= 12'h7F1;
        12'h3B6: sinewave <= 12'h7F1;
        12'h3B7: sinewave <= 12'h7F2;
        12'h3B8: sinewave <= 12'h7F2;
        12'h3B9: sinewave <= 12'h7F2;
        12'h3BA: sinewave <= 12'h7F3;
        12'h3BB: sinewave <= 12'h7F3;
        12'h3BC: sinewave <= 12'h7F3;
        12'h3BD: sinewave <= 12'h7F4;
        12'h3BE: sinewave <= 12'h7F4;
        12'h3BF: sinewave <= 12'h7F4;
        12'h3C0: sinewave <= 12'h7F5;
        12'h3C1: sinewave <= 12'h7F5;
        12'h3C2: sinewave <= 12'h7F5;
        12'h3C3: sinewave <= 12'h7F6;
        12'h3C4: sinewave <= 12'h7F6;
        12'h3C5: sinewave <= 12'h7F6;
        12'h3C6: sinewave <= 12'h7F6;
        12'h3C7: sinewave <= 12'h7F7;
        12'h3C8: sinewave <= 12'h7F7;
        12'h3C9: sinewave <= 12'h7F7;
        12'h3CA: sinewave <= 12'h7F7;
        12'h3CB: sinewave <= 12'h7F8;
        12'h3CC: sinewave <= 12'h7F8;
        12'h3CD: sinewave <= 12'h7F8;
        12'h3CE: sinewave <= 12'h7F8;
        12'h3CF: sinewave <= 12'h7F9;
        12'h3D0: sinewave <= 12'h7F9;
        12'h3D1: sinewave <= 12'h7F9;
        12'h3D2: sinewave <= 12'h7F9;
        12'h3D3: sinewave <= 12'h7FA;
        12'h3D4: sinewave <= 12'h7FA;
        12'h3D5: sinewave <= 12'h7FA;
        12'h3D6: sinewave <= 12'h7FA;
        12'h3D7: sinewave <= 12'h7FA;
        12'h3D8: sinewave <= 12'h7FB;
        12'h3D9: sinewave <= 12'h7FB;
        12'h3DA: sinewave <= 12'h7FB;
        12'h3DB: sinewave <= 12'h7FB;
        12'h3DC: sinewave <= 12'h7FB;
        12'h3DD: sinewave <= 12'h7FC;
        12'h3DE: sinewave <= 12'h7FC;
        12'h3DF: sinewave <= 12'h7FC;
        12'h3E0: sinewave <= 12'h7FC;
        12'h3E1: sinewave <= 12'h7FC;
        12'h3E2: sinewave <= 12'h7FC;
        12'h3E3: sinewave <= 12'h7FC;
        12'h3E4: sinewave <= 12'h7FD;
        12'h3E5: sinewave <= 12'h7FD;
        12'h3E6: sinewave <= 12'h7FD;
        12'h3E7: sinewave <= 12'h7FD;
        12'h3E8: sinewave <= 12'h7FD;
        12'h3E9: sinewave <= 12'h7FD;
        12'h3EA: sinewave <= 12'h7FD;
        12'h3EB: sinewave <= 12'h7FD;
        12'h3EC: sinewave <= 12'h7FE;
        12'h3ED: sinewave <= 12'h7FE;
        12'h3EE: sinewave <= 12'h7FE;
        12'h3EF: sinewave <= 12'h7FE;
        12'h3F0: sinewave <= 12'h7FE;
        12'h3F1: sinewave <= 12'h7FE;
        12'h3F2: sinewave <= 12'h7FE;
        12'h3F3: sinewave <= 12'h7FE;
        12'h3F4: sinewave <= 12'h7FE;
        12'h3F5: sinewave <= 12'h7FE;
        12'h3F6: sinewave <= 12'h7FE;
        12'h3F7: sinewave <= 12'h7FE;
        12'h3F8: sinewave <= 12'h7FE;
        12'h3F9: sinewave <= 12'h7FE;
        12'h3FA: sinewave <= 12'h7FE;
        12'h3FB: sinewave <= 12'h7FE;
        12'h3FC: sinewave <= 12'h7FE;
        12'h3FD: sinewave <= 12'h7FE;
        12'h3FE: sinewave <= 12'h7FE;
        12'h3FF: sinewave <= 12'h7FE;
        12'h400: sinewave <= 12'h7FF;
        12'h401: sinewave <= 12'h7FE;
        12'h402: sinewave <= 12'h7FE;
        12'h403: sinewave <= 12'h7FE;
        12'h404: sinewave <= 12'h7FE;
        12'h405: sinewave <= 12'h7FE;
        12'h406: sinewave <= 12'h7FE;
        12'h407: sinewave <= 12'h7FE;
        12'h408: sinewave <= 12'h7FE;
        12'h409: sinewave <= 12'h7FE;
        12'h40A: sinewave <= 12'h7FE;
        12'h40B: sinewave <= 12'h7FE;
        12'h40C: sinewave <= 12'h7FE;
        12'h40D: sinewave <= 12'h7FE;
        12'h40E: sinewave <= 12'h7FE;
        12'h40F: sinewave <= 12'h7FE;
        12'h410: sinewave <= 12'h7FE;
        12'h411: sinewave <= 12'h7FE;
        12'h412: sinewave <= 12'h7FE;
        12'h413: sinewave <= 12'h7FE;
        12'h414: sinewave <= 12'h7FE;
        12'h415: sinewave <= 12'h7FD;
        12'h416: sinewave <= 12'h7FD;
        12'h417: sinewave <= 12'h7FD;
        12'h418: sinewave <= 12'h7FD;
        12'h419: sinewave <= 12'h7FD;
        12'h41A: sinewave <= 12'h7FD;
        12'h41B: sinewave <= 12'h7FD;
        12'h41C: sinewave <= 12'h7FD;
        12'h41D: sinewave <= 12'h7FC;
        12'h41E: sinewave <= 12'h7FC;
        12'h41F: sinewave <= 12'h7FC;
        12'h420: sinewave <= 12'h7FC;
        12'h421: sinewave <= 12'h7FC;
        12'h422: sinewave <= 12'h7FC;
        12'h423: sinewave <= 12'h7FC;
        12'h424: sinewave <= 12'h7FB;
        12'h425: sinewave <= 12'h7FB;
        12'h426: sinewave <= 12'h7FB;
        12'h427: sinewave <= 12'h7FB;
        12'h428: sinewave <= 12'h7FB;
        12'h429: sinewave <= 12'h7FA;
        12'h42A: sinewave <= 12'h7FA;
        12'h42B: sinewave <= 12'h7FA;
        12'h42C: sinewave <= 12'h7FA;
        12'h42D: sinewave <= 12'h7FA;
        12'h42E: sinewave <= 12'h7F9;
        12'h42F: sinewave <= 12'h7F9;
        12'h430: sinewave <= 12'h7F9;
        12'h431: sinewave <= 12'h7F9;
        12'h432: sinewave <= 12'h7F8;
        12'h433: sinewave <= 12'h7F8;
        12'h434: sinewave <= 12'h7F8;
        12'h435: sinewave <= 12'h7F8;
        12'h436: sinewave <= 12'h7F7;
        12'h437: sinewave <= 12'h7F7;
        12'h438: sinewave <= 12'h7F7;
        12'h439: sinewave <= 12'h7F7;
        12'h43A: sinewave <= 12'h7F6;
        12'h43B: sinewave <= 12'h7F6;
        12'h43C: sinewave <= 12'h7F6;
        12'h43D: sinewave <= 12'h7F6;
        12'h43E: sinewave <= 12'h7F5;
        12'h43F: sinewave <= 12'h7F5;
        12'h440: sinewave <= 12'h7F5;
        12'h441: sinewave <= 12'h7F4;
        12'h442: sinewave <= 12'h7F4;
        12'h443: sinewave <= 12'h7F4;
        12'h444: sinewave <= 12'h7F3;
        12'h445: sinewave <= 12'h7F3;
        12'h446: sinewave <= 12'h7F3;
        12'h447: sinewave <= 12'h7F2;
        12'h448: sinewave <= 12'h7F2;
        12'h449: sinewave <= 12'h7F2;
        12'h44A: sinewave <= 12'h7F1;
        12'h44B: sinewave <= 12'h7F1;
        12'h44C: sinewave <= 12'h7F1;
        12'h44D: sinewave <= 12'h7F0;
        12'h44E: sinewave <= 12'h7F0;
        12'h44F: sinewave <= 12'h7EF;
        12'h450: sinewave <= 12'h7EF;
        12'h451: sinewave <= 12'h7EF;
        12'h452: sinewave <= 12'h7EE;
        12'h453: sinewave <= 12'h7EE;
        12'h454: sinewave <= 12'h7EE;
        12'h455: sinewave <= 12'h7ED;
        12'h456: sinewave <= 12'h7ED;
        12'h457: sinewave <= 12'h7EC;
        12'h458: sinewave <= 12'h7EC;
        12'h459: sinewave <= 12'h7EB;
        12'h45A: sinewave <= 12'h7EB;
        12'h45B: sinewave <= 12'h7EB;
        12'h45C: sinewave <= 12'h7EA;
        12'h45D: sinewave <= 12'h7EA;
        12'h45E: sinewave <= 12'h7E9;
        12'h45F: sinewave <= 12'h7E9;
        12'h460: sinewave <= 12'h7E8;
        12'h461: sinewave <= 12'h7E8;
        12'h462: sinewave <= 12'h7E7;
        12'h463: sinewave <= 12'h7E7;
        12'h464: sinewave <= 12'h7E6;
        12'h465: sinewave <= 12'h7E6;
        12'h466: sinewave <= 12'h7E5;
        12'h467: sinewave <= 12'h7E5;
        12'h468: sinewave <= 12'h7E5;
        12'h469: sinewave <= 12'h7E4;
        12'h46A: sinewave <= 12'h7E3;
        12'h46B: sinewave <= 12'h7E3;
        12'h46C: sinewave <= 12'h7E2;
        12'h46D: sinewave <= 12'h7E2;
        12'h46E: sinewave <= 12'h7E1;
        12'h46F: sinewave <= 12'h7E1;
        12'h470: sinewave <= 12'h7E0;
        12'h471: sinewave <= 12'h7E0;
        12'h472: sinewave <= 12'h7DF;
        12'h473: sinewave <= 12'h7DF;
        12'h474: sinewave <= 12'h7DE;
        12'h475: sinewave <= 12'h7DE;
        12'h476: sinewave <= 12'h7DD;
        12'h477: sinewave <= 12'h7DC;
        12'h478: sinewave <= 12'h7DC;
        12'h479: sinewave <= 12'h7DB;
        12'h47A: sinewave <= 12'h7DB;
        12'h47B: sinewave <= 12'h7DA;
        12'h47C: sinewave <= 12'h7DA;
        12'h47D: sinewave <= 12'h7D9;
        12'h47E: sinewave <= 12'h7D8;
        12'h47F: sinewave <= 12'h7D8;
        12'h480: sinewave <= 12'h7D7;
        12'h481: sinewave <= 12'h7D7;
        12'h482: sinewave <= 12'h7D6;
        12'h483: sinewave <= 12'h7D5;
        12'h484: sinewave <= 12'h7D5;
        12'h485: sinewave <= 12'h7D4;
        12'h486: sinewave <= 12'h7D3;
        12'h487: sinewave <= 12'h7D3;
        12'h488: sinewave <= 12'h7D2;
        12'h489: sinewave <= 12'h7D1;
        12'h48A: sinewave <= 12'h7D1;
        12'h48B: sinewave <= 12'h7D0;
        12'h48C: sinewave <= 12'h7CF;
        12'h48D: sinewave <= 12'h7CF;
        12'h48E: sinewave <= 12'h7CE;
        12'h48F: sinewave <= 12'h7CD;
        12'h490: sinewave <= 12'h7CD;
        12'h491: sinewave <= 12'h7CC;
        12'h492: sinewave <= 12'h7CB;
        12'h493: sinewave <= 12'h7CB;
        12'h494: sinewave <= 12'h7CA;
        12'h495: sinewave <= 12'h7C9;
        12'h496: sinewave <= 12'h7C9;
        12'h497: sinewave <= 12'h7C8;
        12'h498: sinewave <= 12'h7C7;
        12'h499: sinewave <= 12'h7C6;
        12'h49A: sinewave <= 12'h7C6;
        12'h49B: sinewave <= 12'h7C5;
        12'h49C: sinewave <= 12'h7C4;
        12'h49D: sinewave <= 12'h7C3;
        12'h49E: sinewave <= 12'h7C3;
        12'h49F: sinewave <= 12'h7C2;
        12'h4A0: sinewave <= 12'h7C1;
        12'h4A1: sinewave <= 12'h7C0;
        12'h4A2: sinewave <= 12'h7C0;
        12'h4A3: sinewave <= 12'h7BF;
        12'h4A4: sinewave <= 12'h7BE;
        12'h4A5: sinewave <= 12'h7BD;
        12'h4A6: sinewave <= 12'h7BC;
        12'h4A7: sinewave <= 12'h7BC;
        12'h4A8: sinewave <= 12'h7BB;
        12'h4A9: sinewave <= 12'h7BA;
        12'h4AA: sinewave <= 12'h7B9;
        12'h4AB: sinewave <= 12'h7B8;
        12'h4AC: sinewave <= 12'h7B8;
        12'h4AD: sinewave <= 12'h7B7;
        12'h4AE: sinewave <= 12'h7B6;
        12'h4AF: sinewave <= 12'h7B5;
        12'h4B0: sinewave <= 12'h7B4;
        12'h4B1: sinewave <= 12'h7B4;
        12'h4B2: sinewave <= 12'h7B3;
        12'h4B3: sinewave <= 12'h7B2;
        12'h4B4: sinewave <= 12'h7B1;
        12'h4B5: sinewave <= 12'h7B0;
        12'h4B6: sinewave <= 12'h7AF;
        12'h4B7: sinewave <= 12'h7AE;
        12'h4B8: sinewave <= 12'h7AE;
        12'h4B9: sinewave <= 12'h7AD;
        12'h4BA: sinewave <= 12'h7AC;
        12'h4BB: sinewave <= 12'h7AB;
        12'h4BC: sinewave <= 12'h7AA;
        12'h4BD: sinewave <= 12'h7A9;
        12'h4BE: sinewave <= 12'h7A8;
        12'h4BF: sinewave <= 12'h7A7;
        12'h4C0: sinewave <= 12'h7A6;
        12'h4C1: sinewave <= 12'h7A5;
        12'h4C2: sinewave <= 12'h7A5;
        12'h4C3: sinewave <= 12'h7A4;
        12'h4C4: sinewave <= 12'h7A3;
        12'h4C5: sinewave <= 12'h7A2;
        12'h4C6: sinewave <= 12'h7A1;
        12'h4C7: sinewave <= 12'h7A0;
        12'h4C8: sinewave <= 12'h79F;
        12'h4C9: sinewave <= 12'h79E;
        12'h4CA: sinewave <= 12'h79D;
        12'h4CB: sinewave <= 12'h79C;
        12'h4CC: sinewave <= 12'h79B;
        12'h4CD: sinewave <= 12'h79A;
        12'h4CE: sinewave <= 12'h799;
        12'h4CF: sinewave <= 12'h798;
        12'h4D0: sinewave <= 12'h797;
        12'h4D1: sinewave <= 12'h796;
        12'h4D2: sinewave <= 12'h795;
        12'h4D3: sinewave <= 12'h794;
        12'h4D4: sinewave <= 12'h793;
        12'h4D5: sinewave <= 12'h792;
        12'h4D6: sinewave <= 12'h791;
        12'h4D7: sinewave <= 12'h790;
        12'h4D8: sinewave <= 12'h78F;
        12'h4D9: sinewave <= 12'h78E;
        12'h4DA: sinewave <= 12'h78D;
        12'h4DB: sinewave <= 12'h78C;
        12'h4DC: sinewave <= 12'h78B;
        12'h4DD: sinewave <= 12'h78A;
        12'h4DE: sinewave <= 12'h789;
        12'h4DF: sinewave <= 12'h788;
        12'h4E0: sinewave <= 12'h787;
        12'h4E1: sinewave <= 12'h786;
        12'h4E2: sinewave <= 12'h785;
        12'h4E3: sinewave <= 12'h784;
        12'h4E4: sinewave <= 12'h783;
        12'h4E5: sinewave <= 12'h781;
        12'h4E6: sinewave <= 12'h780;
        12'h4E7: sinewave <= 12'h77F;
        12'h4E8: sinewave <= 12'h77E;
        12'h4E9: sinewave <= 12'h77D;
        12'h4EA: sinewave <= 12'h77C;
        12'h4EB: sinewave <= 12'h77B;
        12'h4EC: sinewave <= 12'h77A;
        12'h4ED: sinewave <= 12'h779;
        12'h4EE: sinewave <= 12'h778;
        12'h4EF: sinewave <= 12'h776;
        12'h4F0: sinewave <= 12'h775;
        12'h4F1: sinewave <= 12'h774;
        12'h4F2: sinewave <= 12'h773;
        12'h4F3: sinewave <= 12'h772;
        12'h4F4: sinewave <= 12'h771;
        12'h4F5: sinewave <= 12'h770;
        12'h4F6: sinewave <= 12'h76E;
        12'h4F7: sinewave <= 12'h76D;
        12'h4F8: sinewave <= 12'h76C;
        12'h4F9: sinewave <= 12'h76B;
        12'h4FA: sinewave <= 12'h76A;
        12'h4FB: sinewave <= 12'h769;
        12'h4FC: sinewave <= 12'h767;
        12'h4FD: sinewave <= 12'h766;
        12'h4FE: sinewave <= 12'h765;
        12'h4FF: sinewave <= 12'h764;
        12'h500: sinewave <= 12'h763;
        12'h501: sinewave <= 12'h761;
        12'h502: sinewave <= 12'h760;
        12'h503: sinewave <= 12'h75F;
        12'h504: sinewave <= 12'h75E;
        12'h505: sinewave <= 12'h75D;
        12'h506: sinewave <= 12'h75B;
        12'h507: sinewave <= 12'h75A;
        12'h508: sinewave <= 12'h759;
        12'h509: sinewave <= 12'h758;
        12'h50A: sinewave <= 12'h756;
        12'h50B: sinewave <= 12'h755;
        12'h50C: sinewave <= 12'h754;
        12'h50D: sinewave <= 12'h753;
        12'h50E: sinewave <= 12'h751;
        12'h50F: sinewave <= 12'h750;
        12'h510: sinewave <= 12'h74F;
        12'h511: sinewave <= 12'h74E;
        12'h512: sinewave <= 12'h74C;
        12'h513: sinewave <= 12'h74B;
        12'h514: sinewave <= 12'h74A;
        12'h515: sinewave <= 12'h748;
        12'h516: sinewave <= 12'h747;
        12'h517: sinewave <= 12'h746;
        12'h518: sinewave <= 12'h745;
        12'h519: sinewave <= 12'h743;
        12'h51A: sinewave <= 12'h742;
        12'h51B: sinewave <= 12'h741;
        12'h51C: sinewave <= 12'h73F;
        12'h51D: sinewave <= 12'h73E;
        12'h51E: sinewave <= 12'h73D;
        12'h51F: sinewave <= 12'h73B;
        12'h520: sinewave <= 12'h73A;
        12'h521: sinewave <= 12'h739;
        12'h522: sinewave <= 12'h737;
        12'h523: sinewave <= 12'h736;
        12'h524: sinewave <= 12'h735;
        12'h525: sinewave <= 12'h733;
        12'h526: sinewave <= 12'h732;
        12'h527: sinewave <= 12'h730;
        12'h528: sinewave <= 12'h72F;
        12'h529: sinewave <= 12'h72E;
        12'h52A: sinewave <= 12'h72C;
        12'h52B: sinewave <= 12'h72B;
        12'h52C: sinewave <= 12'h72A;
        12'h52D: sinewave <= 12'h728;
        12'h52E: sinewave <= 12'h727;
        12'h52F: sinewave <= 12'h725;
        12'h530: sinewave <= 12'h724;
        12'h531: sinewave <= 12'h723;
        12'h532: sinewave <= 12'h721;
        12'h533: sinewave <= 12'h720;
        12'h534: sinewave <= 12'h71E;
        12'h535: sinewave <= 12'h71D;
        12'h536: sinewave <= 12'h71B;
        12'h537: sinewave <= 12'h71A;
        12'h538: sinewave <= 12'h718;
        12'h539: sinewave <= 12'h717;
        12'h53A: sinewave <= 12'h716;
        12'h53B: sinewave <= 12'h714;
        12'h53C: sinewave <= 12'h713;
        12'h53D: sinewave <= 12'h711;
        12'h53E: sinewave <= 12'h710;
        12'h53F: sinewave <= 12'h70E;
        12'h540: sinewave <= 12'h70D;
        12'h541: sinewave <= 12'h70B;
        12'h542: sinewave <= 12'h70A;
        12'h543: sinewave <= 12'h708;
        12'h544: sinewave <= 12'h707;
        12'h545: sinewave <= 12'h705;
        12'h546: sinewave <= 12'h704;
        12'h547: sinewave <= 12'h702;
        12'h548: sinewave <= 12'h701;
        12'h549: sinewave <= 12'h6FF;
        12'h54A: sinewave <= 12'h6FE;
        12'h54B: sinewave <= 12'h6FC;
        12'h54C: sinewave <= 12'h6FB;
        12'h54D: sinewave <= 12'h6F9;
        12'h54E: sinewave <= 12'h6F8;
        12'h54F: sinewave <= 12'h6F6;
        12'h550: sinewave <= 12'h6F5;
        12'h551: sinewave <= 12'h6F3;
        12'h552: sinewave <= 12'h6F1;
        12'h553: sinewave <= 12'h6F0;
        12'h554: sinewave <= 12'h6EE;
        12'h555: sinewave <= 12'h6ED;
        12'h556: sinewave <= 12'h6EB;
        12'h557: sinewave <= 12'h6EA;
        12'h558: sinewave <= 12'h6E8;
        12'h559: sinewave <= 12'h6E6;
        12'h55A: sinewave <= 12'h6E5;
        12'h55B: sinewave <= 12'h6E3;
        12'h55C: sinewave <= 12'h6E2;
        12'h55D: sinewave <= 12'h6E0;
        12'h55E: sinewave <= 12'h6DE;
        12'h55F: sinewave <= 12'h6DD;
        12'h560: sinewave <= 12'h6DB;
        12'h561: sinewave <= 12'h6DA;
        12'h562: sinewave <= 12'h6D8;
        12'h563: sinewave <= 12'h6D6;
        12'h564: sinewave <= 12'h6D5;
        12'h565: sinewave <= 12'h6D3;
        12'h566: sinewave <= 12'h6D2;
        12'h567: sinewave <= 12'h6D0;
        12'h568: sinewave <= 12'h6CE;
        12'h569: sinewave <= 12'h6CD;
        12'h56A: sinewave <= 12'h6CB;
        12'h56B: sinewave <= 12'h6C9;
        12'h56C: sinewave <= 12'h6C8;
        12'h56D: sinewave <= 12'h6C6;
        12'h56E: sinewave <= 12'h6C4;
        12'h56F: sinewave <= 12'h6C3;
        12'h570: sinewave <= 12'h6C1;
        12'h571: sinewave <= 12'h6BF;
        12'h572: sinewave <= 12'h6BE;
        12'h573: sinewave <= 12'h6BC;
        12'h574: sinewave <= 12'h6BA;
        12'h575: sinewave <= 12'h6B8;
        12'h576: sinewave <= 12'h6B7;
        12'h577: sinewave <= 12'h6B5;
        12'h578: sinewave <= 12'h6B3;
        12'h579: sinewave <= 12'h6B2;
        12'h57A: sinewave <= 12'h6B0;
        12'h57B: sinewave <= 12'h6AE;
        12'h57C: sinewave <= 12'h6AC;
        12'h57D: sinewave <= 12'h6AB;
        12'h57E: sinewave <= 12'h6A9;
        12'h57F: sinewave <= 12'h6A7;
        12'h580: sinewave <= 12'h6A6;
        12'h581: sinewave <= 12'h6A4;
        12'h582: sinewave <= 12'h6A2;
        12'h583: sinewave <= 12'h6A0;
        12'h584: sinewave <= 12'h69F;
        12'h585: sinewave <= 12'h69D;
        12'h586: sinewave <= 12'h69B;
        12'h587: sinewave <= 12'h699;
        12'h588: sinewave <= 12'h697;
        12'h589: sinewave <= 12'h696;
        12'h58A: sinewave <= 12'h694;
        12'h58B: sinewave <= 12'h692;
        12'h58C: sinewave <= 12'h690;
        12'h58D: sinewave <= 12'h68F;
        12'h58E: sinewave <= 12'h68D;
        12'h58F: sinewave <= 12'h68B;
        12'h590: sinewave <= 12'h689;
        12'h591: sinewave <= 12'h687;
        12'h592: sinewave <= 12'h685;
        12'h593: sinewave <= 12'h684;
        12'h594: sinewave <= 12'h682;
        12'h595: sinewave <= 12'h680;
        12'h596: sinewave <= 12'h67E;
        12'h597: sinewave <= 12'h67C;
        12'h598: sinewave <= 12'h67B;
        12'h599: sinewave <= 12'h679;
        12'h59A: sinewave <= 12'h677;
        12'h59B: sinewave <= 12'h675;
        12'h59C: sinewave <= 12'h673;
        12'h59D: sinewave <= 12'h671;
        12'h59E: sinewave <= 12'h66F;
        12'h59F: sinewave <= 12'h66E;
        12'h5A0: sinewave <= 12'h66C;
        12'h5A1: sinewave <= 12'h66A;
        12'h5A2: sinewave <= 12'h668;
        12'h5A3: sinewave <= 12'h666;
        12'h5A4: sinewave <= 12'h664;
        12'h5A5: sinewave <= 12'h662;
        12'h5A6: sinewave <= 12'h660;
        12'h5A7: sinewave <= 12'h65E;
        12'h5A8: sinewave <= 12'h65D;
        12'h5A9: sinewave <= 12'h65B;
        12'h5AA: sinewave <= 12'h659;
        12'h5AB: sinewave <= 12'h657;
        12'h5AC: sinewave <= 12'h655;
        12'h5AD: sinewave <= 12'h653;
        12'h5AE: sinewave <= 12'h651;
        12'h5AF: sinewave <= 12'h64F;
        12'h5B0: sinewave <= 12'h64D;
        12'h5B1: sinewave <= 12'h64B;
        12'h5B2: sinewave <= 12'h649;
        12'h5B3: sinewave <= 12'h647;
        12'h5B4: sinewave <= 12'h645;
        12'h5B5: sinewave <= 12'h644;
        12'h5B6: sinewave <= 12'h642;
        12'h5B7: sinewave <= 12'h640;
        12'h5B8: sinewave <= 12'h63E;
        12'h5B9: sinewave <= 12'h63C;
        12'h5BA: sinewave <= 12'h63A;
        12'h5BB: sinewave <= 12'h638;
        12'h5BC: sinewave <= 12'h636;
        12'h5BD: sinewave <= 12'h634;
        12'h5BE: sinewave <= 12'h632;
        12'h5BF: sinewave <= 12'h630;
        12'h5C0: sinewave <= 12'h62E;
        12'h5C1: sinewave <= 12'h62C;
        12'h5C2: sinewave <= 12'h62A;
        12'h5C3: sinewave <= 12'h628;
        12'h5C4: sinewave <= 12'h626;
        12'h5C5: sinewave <= 12'h624;
        12'h5C6: sinewave <= 12'h622;
        12'h5C7: sinewave <= 12'h620;
        12'h5C8: sinewave <= 12'h61E;
        12'h5C9: sinewave <= 12'h61C;
        12'h5CA: sinewave <= 12'h61A;
        12'h5CB: sinewave <= 12'h618;
        12'h5CC: sinewave <= 12'h616;
        12'h5CD: sinewave <= 12'h614;
        12'h5CE: sinewave <= 12'h612;
        12'h5CF: sinewave <= 12'h610;
        12'h5D0: sinewave <= 12'h60E;
        12'h5D1: sinewave <= 12'h60B;
        12'h5D2: sinewave <= 12'h609;
        12'h5D3: sinewave <= 12'h607;
        12'h5D4: sinewave <= 12'h605;
        12'h5D5: sinewave <= 12'h603;
        12'h5D6: sinewave <= 12'h601;
        12'h5D7: sinewave <= 12'h5FF;
        12'h5D8: sinewave <= 12'h5FD;
        12'h5D9: sinewave <= 12'h5FB;
        12'h5DA: sinewave <= 12'h5F9;
        12'h5DB: sinewave <= 12'h5F7;
        12'h5DC: sinewave <= 12'h5F5;
        12'h5DD: sinewave <= 12'h5F3;
        12'h5DE: sinewave <= 12'h5F0;
        12'h5DF: sinewave <= 12'h5EE;
        12'h5E0: sinewave <= 12'h5EC;
        12'h5E1: sinewave <= 12'h5EA;
        12'h5E2: sinewave <= 12'h5E8;
        12'h5E3: sinewave <= 12'h5E6;
        12'h5E4: sinewave <= 12'h5E4;
        12'h5E5: sinewave <= 12'h5E2;
        12'h5E6: sinewave <= 12'h5E0;
        12'h5E7: sinewave <= 12'h5DD;
        12'h5E8: sinewave <= 12'h5DB;
        12'h5E9: sinewave <= 12'h5D9;
        12'h5EA: sinewave <= 12'h5D7;
        12'h5EB: sinewave <= 12'h5D5;
        12'h5EC: sinewave <= 12'h5D3;
        12'h5ED: sinewave <= 12'h5D1;
        12'h5EE: sinewave <= 12'h5CE;
        12'h5EF: sinewave <= 12'h5CC;
        12'h5F0: sinewave <= 12'h5CA;
        12'h5F1: sinewave <= 12'h5C8;
        12'h5F2: sinewave <= 12'h5C6;
        12'h5F3: sinewave <= 12'h5C4;
        12'h5F4: sinewave <= 12'h5C1;
        12'h5F5: sinewave <= 12'h5BF;
        12'h5F6: sinewave <= 12'h5BD;
        12'h5F7: sinewave <= 12'h5BB;
        12'h5F8: sinewave <= 12'h5B9;
        12'h5F9: sinewave <= 12'h5B6;
        12'h5FA: sinewave <= 12'h5B4;
        12'h5FB: sinewave <= 12'h5B2;
        12'h5FC: sinewave <= 12'h5B0;
        12'h5FD: sinewave <= 12'h5AE;
        12'h5FE: sinewave <= 12'h5AB;
        12'h5FF: sinewave <= 12'h5A9;
        12'h600: sinewave <= 12'h5A7;
        12'h601: sinewave <= 12'h5A5;
        12'h602: sinewave <= 12'h5A3;
        12'h603: sinewave <= 12'h5A0;
        12'h604: sinewave <= 12'h59E;
        12'h605: sinewave <= 12'h59C;
        12'h606: sinewave <= 12'h59A;
        12'h607: sinewave <= 12'h597;
        12'h608: sinewave <= 12'h595;
        12'h609: sinewave <= 12'h593;
        12'h60A: sinewave <= 12'h591;
        12'h60B: sinewave <= 12'h58E;
        12'h60C: sinewave <= 12'h58C;
        12'h60D: sinewave <= 12'h58A;
        12'h60E: sinewave <= 12'h588;
        12'h60F: sinewave <= 12'h585;
        12'h610: sinewave <= 12'h583;
        12'h611: sinewave <= 12'h581;
        12'h612: sinewave <= 12'h57E;
        12'h613: sinewave <= 12'h57C;
        12'h614: sinewave <= 12'h57A;
        12'h615: sinewave <= 12'h578;
        12'h616: sinewave <= 12'h575;
        12'h617: sinewave <= 12'h573;
        12'h618: sinewave <= 12'h571;
        12'h619: sinewave <= 12'h56E;
        12'h61A: sinewave <= 12'h56C;
        12'h61B: sinewave <= 12'h56A;
        12'h61C: sinewave <= 12'h567;
        12'h61D: sinewave <= 12'h565;
        12'h61E: sinewave <= 12'h563;
        12'h61F: sinewave <= 12'h561;
        12'h620: sinewave <= 12'h55E;
        12'h621: sinewave <= 12'h55C;
        12'h622: sinewave <= 12'h55A;
        12'h623: sinewave <= 12'h557;
        12'h624: sinewave <= 12'h555;
        12'h625: sinewave <= 12'h553;
        12'h626: sinewave <= 12'h550;
        12'h627: sinewave <= 12'h54E;
        12'h628: sinewave <= 12'h54B;
        12'h629: sinewave <= 12'h549;
        12'h62A: sinewave <= 12'h547;
        12'h62B: sinewave <= 12'h544;
        12'h62C: sinewave <= 12'h542;
        12'h62D: sinewave <= 12'h540;
        12'h62E: sinewave <= 12'h53D;
        12'h62F: sinewave <= 12'h53B;
        12'h630: sinewave <= 12'h539;
        12'h631: sinewave <= 12'h536;
        12'h632: sinewave <= 12'h534;
        12'h633: sinewave <= 12'h531;
        12'h634: sinewave <= 12'h52F;
        12'h635: sinewave <= 12'h52D;
        12'h636: sinewave <= 12'h52A;
        12'h637: sinewave <= 12'h528;
        12'h638: sinewave <= 12'h525;
        12'h639: sinewave <= 12'h523;
        12'h63A: sinewave <= 12'h521;
        12'h63B: sinewave <= 12'h51E;
        12'h63C: sinewave <= 12'h51C;
        12'h63D: sinewave <= 12'h519;
        12'h63E: sinewave <= 12'h517;
        12'h63F: sinewave <= 12'h515;
        12'h640: sinewave <= 12'h512;
        12'h641: sinewave <= 12'h510;
        12'h642: sinewave <= 12'h50D;
        12'h643: sinewave <= 12'h50B;
        12'h644: sinewave <= 12'h508;
        12'h645: sinewave <= 12'h506;
        12'h646: sinewave <= 12'h503;
        12'h647: sinewave <= 12'h501;
        12'h648: sinewave <= 12'h4FF;
        12'h649: sinewave <= 12'h4FC;
        12'h64A: sinewave <= 12'h4FA;
        12'h64B: sinewave <= 12'h4F7;
        12'h64C: sinewave <= 12'h4F5;
        12'h64D: sinewave <= 12'h4F2;
        12'h64E: sinewave <= 12'h4F0;
        12'h64F: sinewave <= 12'h4ED;
        12'h650: sinewave <= 12'h4EB;
        12'h651: sinewave <= 12'h4E8;
        12'h652: sinewave <= 12'h4E6;
        12'h653: sinewave <= 12'h4E3;
        12'h654: sinewave <= 12'h4E1;
        12'h655: sinewave <= 12'h4DE;
        12'h656: sinewave <= 12'h4DC;
        12'h657: sinewave <= 12'h4D9;
        12'h658: sinewave <= 12'h4D7;
        12'h659: sinewave <= 12'h4D4;
        12'h65A: sinewave <= 12'h4D2;
        12'h65B: sinewave <= 12'h4CF;
        12'h65C: sinewave <= 12'h4CD;
        12'h65D: sinewave <= 12'h4CA;
        12'h65E: sinewave <= 12'h4C8;
        12'h65F: sinewave <= 12'h4C5;
        12'h660: sinewave <= 12'h4C3;
        12'h661: sinewave <= 12'h4C0;
        12'h662: sinewave <= 12'h4BE;
        12'h663: sinewave <= 12'h4BB;
        12'h664: sinewave <= 12'h4B9;
        12'h665: sinewave <= 12'h4B6;
        12'h666: sinewave <= 12'h4B4;
        12'h667: sinewave <= 12'h4B1;
        12'h668: sinewave <= 12'h4AF;
        12'h669: sinewave <= 12'h4AC;
        12'h66A: sinewave <= 12'h4AA;
        12'h66B: sinewave <= 12'h4A7;
        12'h66C: sinewave <= 12'h4A4;
        12'h66D: sinewave <= 12'h4A2;
        12'h66E: sinewave <= 12'h49F;
        12'h66F: sinewave <= 12'h49D;
        12'h670: sinewave <= 12'h49A;
        12'h671: sinewave <= 12'h498;
        12'h672: sinewave <= 12'h495;
        12'h673: sinewave <= 12'h492;
        12'h674: sinewave <= 12'h490;
        12'h675: sinewave <= 12'h48D;
        12'h676: sinewave <= 12'h48B;
        12'h677: sinewave <= 12'h488;
        12'h678: sinewave <= 12'h486;
        12'h679: sinewave <= 12'h483;
        12'h67A: sinewave <= 12'h480;
        12'h67B: sinewave <= 12'h47E;
        12'h67C: sinewave <= 12'h47B;
        12'h67D: sinewave <= 12'h479;
        12'h67E: sinewave <= 12'h476;
        12'h67F: sinewave <= 12'h473;
        12'h680: sinewave <= 12'h471;
        12'h681: sinewave <= 12'h46E;
        12'h682: sinewave <= 12'h46C;
        12'h683: sinewave <= 12'h469;
        12'h684: sinewave <= 12'h466;
        12'h685: sinewave <= 12'h464;
        12'h686: sinewave <= 12'h461;
        12'h687: sinewave <= 12'h45E;
        12'h688: sinewave <= 12'h45C;
        12'h689: sinewave <= 12'h459;
        12'h68A: sinewave <= 12'h457;
        12'h68B: sinewave <= 12'h454;
        12'h68C: sinewave <= 12'h451;
        12'h68D: sinewave <= 12'h44F;
        12'h68E: sinewave <= 12'h44C;
        12'h68F: sinewave <= 12'h449;
        12'h690: sinewave <= 12'h447;
        12'h691: sinewave <= 12'h444;
        12'h692: sinewave <= 12'h441;
        12'h693: sinewave <= 12'h43F;
        12'h694: sinewave <= 12'h43C;
        12'h695: sinewave <= 12'h439;
        12'h696: sinewave <= 12'h437;
        12'h697: sinewave <= 12'h434;
        12'h698: sinewave <= 12'h431;
        12'h699: sinewave <= 12'h42F;
        12'h69A: sinewave <= 12'h42C;
        12'h69B: sinewave <= 12'h429;
        12'h69C: sinewave <= 12'h427;
        12'h69D: sinewave <= 12'h424;
        12'h69E: sinewave <= 12'h421;
        12'h69F: sinewave <= 12'h41F;
        12'h6A0: sinewave <= 12'h41C;
        12'h6A1: sinewave <= 12'h419;
        12'h6A2: sinewave <= 12'h416;
        12'h6A3: sinewave <= 12'h414;
        12'h6A4: sinewave <= 12'h411;
        12'h6A5: sinewave <= 12'h40E;
        12'h6A6: sinewave <= 12'h40C;
        12'h6A7: sinewave <= 12'h409;
        12'h6A8: sinewave <= 12'h406;
        12'h6A9: sinewave <= 12'h404;
        12'h6AA: sinewave <= 12'h401;
        12'h6AB: sinewave <= 12'h3FE;
        12'h6AC: sinewave <= 12'h3FB;
        12'h6AD: sinewave <= 12'h3F9;
        12'h6AE: sinewave <= 12'h3F6;
        12'h6AF: sinewave <= 12'h3F3;
        12'h6B0: sinewave <= 12'h3F0;
        12'h6B1: sinewave <= 12'h3EE;
        12'h6B2: sinewave <= 12'h3EB;
        12'h6B3: sinewave <= 12'h3E8;
        12'h6B4: sinewave <= 12'h3E6;
        12'h6B5: sinewave <= 12'h3E3;
        12'h6B6: sinewave <= 12'h3E0;
        12'h6B7: sinewave <= 12'h3DD;
        12'h6B8: sinewave <= 12'h3DB;
        12'h6B9: sinewave <= 12'h3D8;
        12'h6BA: sinewave <= 12'h3D5;
        12'h6BB: sinewave <= 12'h3D2;
        12'h6BC: sinewave <= 12'h3D0;
        12'h6BD: sinewave <= 12'h3CD;
        12'h6BE: sinewave <= 12'h3CA;
        12'h6BF: sinewave <= 12'h3C7;
        12'h6C0: sinewave <= 12'h3C4;
        12'h6C1: sinewave <= 12'h3C2;
        12'h6C2: sinewave <= 12'h3BF;
        12'h6C3: sinewave <= 12'h3BC;
        12'h6C4: sinewave <= 12'h3B9;
        12'h6C5: sinewave <= 12'h3B7;
        12'h6C6: sinewave <= 12'h3B4;
        12'h6C7: sinewave <= 12'h3B1;
        12'h6C8: sinewave <= 12'h3AE;
        12'h6C9: sinewave <= 12'h3AB;
        12'h6CA: sinewave <= 12'h3A9;
        12'h6CB: sinewave <= 12'h3A6;
        12'h6CC: sinewave <= 12'h3A3;
        12'h6CD: sinewave <= 12'h3A0;
        12'h6CE: sinewave <= 12'h39D;
        12'h6CF: sinewave <= 12'h39B;
        12'h6D0: sinewave <= 12'h398;
        12'h6D1: sinewave <= 12'h395;
        12'h6D2: sinewave <= 12'h392;
        12'h6D3: sinewave <= 12'h38F;
        12'h6D4: sinewave <= 12'h38D;
        12'h6D5: sinewave <= 12'h38A;
        12'h6D6: sinewave <= 12'h387;
        12'h6D7: sinewave <= 12'h384;
        12'h6D8: sinewave <= 12'h381;
        12'h6D9: sinewave <= 12'h37F;
        12'h6DA: sinewave <= 12'h37C;
        12'h6DB: sinewave <= 12'h379;
        12'h6DC: sinewave <= 12'h376;
        12'h6DD: sinewave <= 12'h373;
        12'h6DE: sinewave <= 12'h370;
        12'h6DF: sinewave <= 12'h36E;
        12'h6E0: sinewave <= 12'h36B;
        12'h6E1: sinewave <= 12'h368;
        12'h6E2: sinewave <= 12'h365;
        12'h6E3: sinewave <= 12'h362;
        12'h6E4: sinewave <= 12'h35F;
        12'h6E5: sinewave <= 12'h35C;
        12'h6E6: sinewave <= 12'h35A;
        12'h6E7: sinewave <= 12'h357;
        12'h6E8: sinewave <= 12'h354;
        12'h6E9: sinewave <= 12'h351;
        12'h6EA: sinewave <= 12'h34E;
        12'h6EB: sinewave <= 12'h34B;
        12'h6EC: sinewave <= 12'h348;
        12'h6ED: sinewave <= 12'h346;
        12'h6EE: sinewave <= 12'h343;
        12'h6EF: sinewave <= 12'h340;
        12'h6F0: sinewave <= 12'h33D;
        12'h6F1: sinewave <= 12'h33A;
        12'h6F2: sinewave <= 12'h337;
        12'h6F3: sinewave <= 12'h334;
        12'h6F4: sinewave <= 12'h332;
        12'h6F5: sinewave <= 12'h32F;
        12'h6F6: sinewave <= 12'h32C;
        12'h6F7: sinewave <= 12'h329;
        12'h6F8: sinewave <= 12'h326;
        12'h6F9: sinewave <= 12'h323;
        12'h6FA: sinewave <= 12'h320;
        12'h6FB: sinewave <= 12'h31D;
        12'h6FC: sinewave <= 12'h31A;
        12'h6FD: sinewave <= 12'h318;
        12'h6FE: sinewave <= 12'h315;
        12'h6FF: sinewave <= 12'h312;
        12'h700: sinewave <= 12'h30F;
        12'h701: sinewave <= 12'h30C;
        12'h702: sinewave <= 12'h309;
        12'h703: sinewave <= 12'h306;
        12'h704: sinewave <= 12'h303;
        12'h705: sinewave <= 12'h300;
        12'h706: sinewave <= 12'h2FD;
        12'h707: sinewave <= 12'h2FB;
        12'h708: sinewave <= 12'h2F8;
        12'h709: sinewave <= 12'h2F5;
        12'h70A: sinewave <= 12'h2F2;
        12'h70B: sinewave <= 12'h2EF;
        12'h70C: sinewave <= 12'h2EC;
        12'h70D: sinewave <= 12'h2E9;
        12'h70E: sinewave <= 12'h2E6;
        12'h70F: sinewave <= 12'h2E3;
        12'h710: sinewave <= 12'h2E0;
        12'h711: sinewave <= 12'h2DD;
        12'h712: sinewave <= 12'h2DA;
        12'h713: sinewave <= 12'h2D7;
        12'h714: sinewave <= 12'h2D4;
        12'h715: sinewave <= 12'h2D2;
        12'h716: sinewave <= 12'h2CF;
        12'h717: sinewave <= 12'h2CC;
        12'h718: sinewave <= 12'h2C9;
        12'h719: sinewave <= 12'h2C6;
        12'h71A: sinewave <= 12'h2C3;
        12'h71B: sinewave <= 12'h2C0;
        12'h71C: sinewave <= 12'h2BD;
        12'h71D: sinewave <= 12'h2BA;
        12'h71E: sinewave <= 12'h2B7;
        12'h71F: sinewave <= 12'h2B4;
        12'h720: sinewave <= 12'h2B1;
        12'h721: sinewave <= 12'h2AE;
        12'h722: sinewave <= 12'h2AB;
        12'h723: sinewave <= 12'h2A8;
        12'h724: sinewave <= 12'h2A5;
        12'h725: sinewave <= 12'h2A2;
        12'h726: sinewave <= 12'h29F;
        12'h727: sinewave <= 12'h29C;
        12'h728: sinewave <= 12'h299;
        12'h729: sinewave <= 12'h296;
        12'h72A: sinewave <= 12'h293;
        12'h72B: sinewave <= 12'h290;
        12'h72C: sinewave <= 12'h28E;
        12'h72D: sinewave <= 12'h28B;
        12'h72E: sinewave <= 12'h288;
        12'h72F: sinewave <= 12'h285;
        12'h730: sinewave <= 12'h282;
        12'h731: sinewave <= 12'h27F;
        12'h732: sinewave <= 12'h27C;
        12'h733: sinewave <= 12'h279;
        12'h734: sinewave <= 12'h276;
        12'h735: sinewave <= 12'h273;
        12'h736: sinewave <= 12'h270;
        12'h737: sinewave <= 12'h26D;
        12'h738: sinewave <= 12'h26A;
        12'h739: sinewave <= 12'h267;
        12'h73A: sinewave <= 12'h264;
        12'h73B: sinewave <= 12'h261;
        12'h73C: sinewave <= 12'h25E;
        12'h73D: sinewave <= 12'h25B;
        12'h73E: sinewave <= 12'h258;
        12'h73F: sinewave <= 12'h255;
        12'h740: sinewave <= 12'h252;
        12'h741: sinewave <= 12'h24F;
        12'h742: sinewave <= 12'h24C;
        12'h743: sinewave <= 12'h249;
        12'h744: sinewave <= 12'h246;
        12'h745: sinewave <= 12'h243;
        12'h746: sinewave <= 12'h240;
        12'h747: sinewave <= 12'h23D;
        12'h748: sinewave <= 12'h23A;
        12'h749: sinewave <= 12'h237;
        12'h74A: sinewave <= 12'h234;
        12'h74B: sinewave <= 12'h231;
        12'h74C: sinewave <= 12'h22E;
        12'h74D: sinewave <= 12'h22B;
        12'h74E: sinewave <= 12'h228;
        12'h74F: sinewave <= 12'h224;
        12'h750: sinewave <= 12'h221;
        12'h751: sinewave <= 12'h21E;
        12'h752: sinewave <= 12'h21B;
        12'h753: sinewave <= 12'h218;
        12'h754: sinewave <= 12'h215;
        12'h755: sinewave <= 12'h212;
        12'h756: sinewave <= 12'h20F;
        12'h757: sinewave <= 12'h20C;
        12'h758: sinewave <= 12'h209;
        12'h759: sinewave <= 12'h206;
        12'h75A: sinewave <= 12'h203;
        12'h75B: sinewave <= 12'h200;
        12'h75C: sinewave <= 12'h1FD;
        12'h75D: sinewave <= 12'h1FA;
        12'h75E: sinewave <= 12'h1F7;
        12'h75F: sinewave <= 12'h1F4;
        12'h760: sinewave <= 12'h1F1;
        12'h761: sinewave <= 12'h1EE;
        12'h762: sinewave <= 12'h1EB;
        12'h763: sinewave <= 12'h1E8;
        12'h764: sinewave <= 12'h1E5;
        12'h765: sinewave <= 12'h1E2;
        12'h766: sinewave <= 12'h1DF;
        12'h767: sinewave <= 12'h1DC;
        12'h768: sinewave <= 12'h1D8;
        12'h769: sinewave <= 12'h1D5;
        12'h76A: sinewave <= 12'h1D2;
        12'h76B: sinewave <= 12'h1CF;
        12'h76C: sinewave <= 12'h1CC;
        12'h76D: sinewave <= 12'h1C9;
        12'h76E: sinewave <= 12'h1C6;
        12'h76F: sinewave <= 12'h1C3;
        12'h770: sinewave <= 12'h1C0;
        12'h771: sinewave <= 12'h1BD;
        12'h772: sinewave <= 12'h1BA;
        12'h773: sinewave <= 12'h1B7;
        12'h774: sinewave <= 12'h1B4;
        12'h775: sinewave <= 12'h1B1;
        12'h776: sinewave <= 12'h1AE;
        12'h777: sinewave <= 12'h1AB;
        12'h778: sinewave <= 12'h1A7;
        12'h779: sinewave <= 12'h1A4;
        12'h77A: sinewave <= 12'h1A1;
        12'h77B: sinewave <= 12'h19E;
        12'h77C: sinewave <= 12'h19B;
        12'h77D: sinewave <= 12'h198;
        12'h77E: sinewave <= 12'h195;
        12'h77F: sinewave <= 12'h192;
        12'h780: sinewave <= 12'h18F;
        12'h781: sinewave <= 12'h18C;
        12'h782: sinewave <= 12'h189;
        12'h783: sinewave <= 12'h186;
        12'h784: sinewave <= 12'h183;
        12'h785: sinewave <= 12'h17F;
        12'h786: sinewave <= 12'h17C;
        12'h787: sinewave <= 12'h179;
        12'h788: sinewave <= 12'h176;
        12'h789: sinewave <= 12'h173;
        12'h78A: sinewave <= 12'h170;
        12'h78B: sinewave <= 12'h16D;
        12'h78C: sinewave <= 12'h16A;
        12'h78D: sinewave <= 12'h167;
        12'h78E: sinewave <= 12'h164;
        12'h78F: sinewave <= 12'h161;
        12'h790: sinewave <= 12'h15D;
        12'h791: sinewave <= 12'h15A;
        12'h792: sinewave <= 12'h157;
        12'h793: sinewave <= 12'h154;
        12'h794: sinewave <= 12'h151;
        12'h795: sinewave <= 12'h14E;
        12'h796: sinewave <= 12'h14B;
        12'h797: sinewave <= 12'h148;
        12'h798: sinewave <= 12'h145;
        12'h799: sinewave <= 12'h142;
        12'h79A: sinewave <= 12'h13E;
        12'h79B: sinewave <= 12'h13B;
        12'h79C: sinewave <= 12'h138;
        12'h79D: sinewave <= 12'h135;
        12'h79E: sinewave <= 12'h132;
        12'h79F: sinewave <= 12'h12F;
        12'h7A0: sinewave <= 12'h12C;
        12'h7A1: sinewave <= 12'h129;
        12'h7A2: sinewave <= 12'h126;
        12'h7A3: sinewave <= 12'h123;
        12'h7A4: sinewave <= 12'h11F;
        12'h7A5: sinewave <= 12'h11C;
        12'h7A6: sinewave <= 12'h119;
        12'h7A7: sinewave <= 12'h116;
        12'h7A8: sinewave <= 12'h113;
        12'h7A9: sinewave <= 12'h110;
        12'h7AA: sinewave <= 12'h10D;
        12'h7AB: sinewave <= 12'h10A;
        12'h7AC: sinewave <= 12'h107;
        12'h7AD: sinewave <= 12'h103;
        12'h7AE: sinewave <= 12'h100;
        12'h7AF: sinewave <= 12'h0FD;
        12'h7B0: sinewave <= 12'h0FA;
        12'h7B1: sinewave <= 12'h0F7;
        12'h7B2: sinewave <= 12'h0F4;
        12'h7B3: sinewave <= 12'h0F1;
        12'h7B4: sinewave <= 12'h0EE;
        12'h7B5: sinewave <= 12'h0EA;
        12'h7B6: sinewave <= 12'h0E7;
        12'h7B7: sinewave <= 12'h0E4;
        12'h7B8: sinewave <= 12'h0E1;
        12'h7B9: sinewave <= 12'h0DE;
        12'h7BA: sinewave <= 12'h0DB;
        12'h7BB: sinewave <= 12'h0D8;
        12'h7BC: sinewave <= 12'h0D5;
        12'h7BD: sinewave <= 12'h0D2;
        12'h7BE: sinewave <= 12'h0CE;
        12'h7BF: sinewave <= 12'h0CB;
        12'h7C0: sinewave <= 12'h0C8;
        12'h7C1: sinewave <= 12'h0C5;
        12'h7C2: sinewave <= 12'h0C2;
        12'h7C3: sinewave <= 12'h0BF;
        12'h7C4: sinewave <= 12'h0BC;
        12'h7C5: sinewave <= 12'h0B9;
        12'h7C6: sinewave <= 12'h0B5;
        12'h7C7: sinewave <= 12'h0B2;
        12'h7C8: sinewave <= 12'h0AF;
        12'h7C9: sinewave <= 12'h0AC;
        12'h7CA: sinewave <= 12'h0A9;
        12'h7CB: sinewave <= 12'h0A6;
        12'h7CC: sinewave <= 12'h0A3;
        12'h7CD: sinewave <= 12'h09F;
        12'h7CE: sinewave <= 12'h09C;
        12'h7CF: sinewave <= 12'h099;
        12'h7D0: sinewave <= 12'h096;
        12'h7D1: sinewave <= 12'h093;
        12'h7D2: sinewave <= 12'h090;
        12'h7D3: sinewave <= 12'h08D;
        12'h7D4: sinewave <= 12'h08A;
        12'h7D5: sinewave <= 12'h086;
        12'h7D6: sinewave <= 12'h083;
        12'h7D7: sinewave <= 12'h080;
        12'h7D8: sinewave <= 12'h07D;
        12'h7D9: sinewave <= 12'h07A;
        12'h7DA: sinewave <= 12'h077;
        12'h7DB: sinewave <= 12'h074;
        12'h7DC: sinewave <= 12'h070;
        12'h7DD: sinewave <= 12'h06D;
        12'h7DE: sinewave <= 12'h06A;
        12'h7DF: sinewave <= 12'h067;
        12'h7E0: sinewave <= 12'h064;
        12'h7E1: sinewave <= 12'h061;
        12'h7E2: sinewave <= 12'h05E;
        12'h7E3: sinewave <= 12'h05B;
        12'h7E4: sinewave <= 12'h057;
        12'h7E5: sinewave <= 12'h054;
        12'h7E6: sinewave <= 12'h051;
        12'h7E7: sinewave <= 12'h04E;
        12'h7E8: sinewave <= 12'h04B;
        12'h7E9: sinewave <= 12'h048;
        12'h7EA: sinewave <= 12'h045;
        12'h7EB: sinewave <= 12'h041;
        12'h7EC: sinewave <= 12'h03E;
        12'h7ED: sinewave <= 12'h03B;
        12'h7EE: sinewave <= 12'h038;
        12'h7EF: sinewave <= 12'h035;
        12'h7F0: sinewave <= 12'h032;
        12'h7F1: sinewave <= 12'h02F;
        12'h7F2: sinewave <= 12'h02B;
        12'h7F3: sinewave <= 12'h028;
        12'h7F4: sinewave <= 12'h025;
        12'h7F5: sinewave <= 12'h022;
        12'h7F6: sinewave <= 12'h01F;
        12'h7F7: sinewave <= 12'h01C;
        12'h7F8: sinewave <= 12'h019;
        12'h7F9: sinewave <= 12'h015;
        12'h7FA: sinewave <= 12'h012;
        12'h7FB: sinewave <= 12'h00F;
        12'h7FC: sinewave <= 12'h00C;
        12'h7FD: sinewave <= 12'h009;
        12'h7FE: sinewave <= 12'h006;
        12'h7FF: sinewave <= 12'h003;
        12'h800: sinewave <= 12'h000;
        12'h801: sinewave <= 12'hFFD;
        12'h802: sinewave <= 12'hFFA;
        12'h803: sinewave <= 12'hFF7;
        12'h804: sinewave <= 12'hFF4;
        12'h805: sinewave <= 12'hFF1;
        12'h806: sinewave <= 12'hFEE;
        12'h807: sinewave <= 12'hFEB;
        12'h808: sinewave <= 12'hFE7;
        12'h809: sinewave <= 12'hFE4;
        12'h80A: sinewave <= 12'hFE1;
        12'h80B: sinewave <= 12'hFDE;
        12'h80C: sinewave <= 12'hFDB;
        12'h80D: sinewave <= 12'hFD8;
        12'h80E: sinewave <= 12'hFD5;
        12'h80F: sinewave <= 12'hFD1;
        12'h810: sinewave <= 12'hFCE;
        12'h811: sinewave <= 12'hFCB;
        12'h812: sinewave <= 12'hFC8;
        12'h813: sinewave <= 12'hFC5;
        12'h814: sinewave <= 12'hFC2;
        12'h815: sinewave <= 12'hFBF;
        12'h816: sinewave <= 12'hFBB;
        12'h817: sinewave <= 12'hFB8;
        12'h818: sinewave <= 12'hFB5;
        12'h819: sinewave <= 12'hFB2;
        12'h81A: sinewave <= 12'hFAF;
        12'h81B: sinewave <= 12'hFAC;
        12'h81C: sinewave <= 12'hFA9;
        12'h81D: sinewave <= 12'hFA5;
        12'h81E: sinewave <= 12'hFA2;
        12'h81F: sinewave <= 12'hF9F;
        12'h820: sinewave <= 12'hF9C;
        12'h821: sinewave <= 12'hF99;
        12'h822: sinewave <= 12'hF96;
        12'h823: sinewave <= 12'hF93;
        12'h824: sinewave <= 12'hF90;
        12'h825: sinewave <= 12'hF8C;
        12'h826: sinewave <= 12'hF89;
        12'h827: sinewave <= 12'hF86;
        12'h828: sinewave <= 12'hF83;
        12'h829: sinewave <= 12'hF80;
        12'h82A: sinewave <= 12'hF7D;
        12'h82B: sinewave <= 12'hF7A;
        12'h82C: sinewave <= 12'hF76;
        12'h82D: sinewave <= 12'hF73;
        12'h82E: sinewave <= 12'hF70;
        12'h82F: sinewave <= 12'hF6D;
        12'h830: sinewave <= 12'hF6A;
        12'h831: sinewave <= 12'hF67;
        12'h832: sinewave <= 12'hF64;
        12'h833: sinewave <= 12'hF61;
        12'h834: sinewave <= 12'hF5D;
        12'h835: sinewave <= 12'hF5A;
        12'h836: sinewave <= 12'hF57;
        12'h837: sinewave <= 12'hF54;
        12'h838: sinewave <= 12'hF51;
        12'h839: sinewave <= 12'hF4E;
        12'h83A: sinewave <= 12'hF4B;
        12'h83B: sinewave <= 12'hF47;
        12'h83C: sinewave <= 12'hF44;
        12'h83D: sinewave <= 12'hF41;
        12'h83E: sinewave <= 12'hF3E;
        12'h83F: sinewave <= 12'hF3B;
        12'h840: sinewave <= 12'hF38;
        12'h841: sinewave <= 12'hF35;
        12'h842: sinewave <= 12'hF32;
        12'h843: sinewave <= 12'hF2E;
        12'h844: sinewave <= 12'hF2B;
        12'h845: sinewave <= 12'hF28;
        12'h846: sinewave <= 12'hF25;
        12'h847: sinewave <= 12'hF22;
        12'h848: sinewave <= 12'hF1F;
        12'h849: sinewave <= 12'hF1C;
        12'h84A: sinewave <= 12'hF19;
        12'h84B: sinewave <= 12'hF16;
        12'h84C: sinewave <= 12'hF12;
        12'h84D: sinewave <= 12'hF0F;
        12'h84E: sinewave <= 12'hF0C;
        12'h84F: sinewave <= 12'hF09;
        12'h850: sinewave <= 12'hF06;
        12'h851: sinewave <= 12'hF03;
        12'h852: sinewave <= 12'hF00;
        12'h853: sinewave <= 12'hEFD;
        12'h854: sinewave <= 12'hEF9;
        12'h855: sinewave <= 12'hEF6;
        12'h856: sinewave <= 12'hEF3;
        12'h857: sinewave <= 12'hEF0;
        12'h858: sinewave <= 12'hEED;
        12'h859: sinewave <= 12'hEEA;
        12'h85A: sinewave <= 12'hEE7;
        12'h85B: sinewave <= 12'hEE4;
        12'h85C: sinewave <= 12'hEE1;
        12'h85D: sinewave <= 12'hEDD;
        12'h85E: sinewave <= 12'hEDA;
        12'h85F: sinewave <= 12'hED7;
        12'h860: sinewave <= 12'hED4;
        12'h861: sinewave <= 12'hED1;
        12'h862: sinewave <= 12'hECE;
        12'h863: sinewave <= 12'hECB;
        12'h864: sinewave <= 12'hEC8;
        12'h865: sinewave <= 12'hEC5;
        12'h866: sinewave <= 12'hEC2;
        12'h867: sinewave <= 12'hEBE;
        12'h868: sinewave <= 12'hEBB;
        12'h869: sinewave <= 12'hEB8;
        12'h86A: sinewave <= 12'hEB5;
        12'h86B: sinewave <= 12'hEB2;
        12'h86C: sinewave <= 12'hEAF;
        12'h86D: sinewave <= 12'hEAC;
        12'h86E: sinewave <= 12'hEA9;
        12'h86F: sinewave <= 12'hEA6;
        12'h870: sinewave <= 12'hEA3;
        12'h871: sinewave <= 12'hE9F;
        12'h872: sinewave <= 12'hE9C;
        12'h873: sinewave <= 12'hE99;
        12'h874: sinewave <= 12'hE96;
        12'h875: sinewave <= 12'hE93;
        12'h876: sinewave <= 12'hE90;
        12'h877: sinewave <= 12'hE8D;
        12'h878: sinewave <= 12'hE8A;
        12'h879: sinewave <= 12'hE87;
        12'h87A: sinewave <= 12'hE84;
        12'h87B: sinewave <= 12'hE81;
        12'h87C: sinewave <= 12'hE7D;
        12'h87D: sinewave <= 12'hE7A;
        12'h87E: sinewave <= 12'hE77;
        12'h87F: sinewave <= 12'hE74;
        12'h880: sinewave <= 12'hE71;
        12'h881: sinewave <= 12'hE6E;
        12'h882: sinewave <= 12'hE6B;
        12'h883: sinewave <= 12'hE68;
        12'h884: sinewave <= 12'hE65;
        12'h885: sinewave <= 12'hE62;
        12'h886: sinewave <= 12'hE5F;
        12'h887: sinewave <= 12'hE5C;
        12'h888: sinewave <= 12'hE59;
        12'h889: sinewave <= 12'hE55;
        12'h88A: sinewave <= 12'hE52;
        12'h88B: sinewave <= 12'hE4F;
        12'h88C: sinewave <= 12'hE4C;
        12'h88D: sinewave <= 12'hE49;
        12'h88E: sinewave <= 12'hE46;
        12'h88F: sinewave <= 12'hE43;
        12'h890: sinewave <= 12'hE40;
        12'h891: sinewave <= 12'hE3D;
        12'h892: sinewave <= 12'hE3A;
        12'h893: sinewave <= 12'hE37;
        12'h894: sinewave <= 12'hE34;
        12'h895: sinewave <= 12'hE31;
        12'h896: sinewave <= 12'hE2E;
        12'h897: sinewave <= 12'hE2B;
        12'h898: sinewave <= 12'hE28;
        12'h899: sinewave <= 12'hE24;
        12'h89A: sinewave <= 12'hE21;
        12'h89B: sinewave <= 12'hE1E;
        12'h89C: sinewave <= 12'hE1B;
        12'h89D: sinewave <= 12'hE18;
        12'h89E: sinewave <= 12'hE15;
        12'h89F: sinewave <= 12'hE12;
        12'h8A0: sinewave <= 12'hE0F;
        12'h8A1: sinewave <= 12'hE0C;
        12'h8A2: sinewave <= 12'hE09;
        12'h8A3: sinewave <= 12'hE06;
        12'h8A4: sinewave <= 12'hE03;
        12'h8A5: sinewave <= 12'hE00;
        12'h8A6: sinewave <= 12'hDFD;
        12'h8A7: sinewave <= 12'hDFA;
        12'h8A8: sinewave <= 12'hDF7;
        12'h8A9: sinewave <= 12'hDF4;
        12'h8AA: sinewave <= 12'hDF1;
        12'h8AB: sinewave <= 12'hDEE;
        12'h8AC: sinewave <= 12'hDEB;
        12'h8AD: sinewave <= 12'hDE8;
        12'h8AE: sinewave <= 12'hDE5;
        12'h8AF: sinewave <= 12'hDE2;
        12'h8B0: sinewave <= 12'hDDF;
        12'h8B1: sinewave <= 12'hDDC;
        12'h8B2: sinewave <= 12'hDD8;
        12'h8B3: sinewave <= 12'hDD5;
        12'h8B4: sinewave <= 12'hDD2;
        12'h8B5: sinewave <= 12'hDCF;
        12'h8B6: sinewave <= 12'hDCC;
        12'h8B7: sinewave <= 12'hDC9;
        12'h8B8: sinewave <= 12'hDC6;
        12'h8B9: sinewave <= 12'hDC3;
        12'h8BA: sinewave <= 12'hDC0;
        12'h8BB: sinewave <= 12'hDBD;
        12'h8BC: sinewave <= 12'hDBA;
        12'h8BD: sinewave <= 12'hDB7;
        12'h8BE: sinewave <= 12'hDB4;
        12'h8BF: sinewave <= 12'hDB1;
        12'h8C0: sinewave <= 12'hDAE;
        12'h8C1: sinewave <= 12'hDAB;
        12'h8C2: sinewave <= 12'hDA8;
        12'h8C3: sinewave <= 12'hDA5;
        12'h8C4: sinewave <= 12'hDA2;
        12'h8C5: sinewave <= 12'hD9F;
        12'h8C6: sinewave <= 12'hD9C;
        12'h8C7: sinewave <= 12'hD99;
        12'h8C8: sinewave <= 12'hD96;
        12'h8C9: sinewave <= 12'hD93;
        12'h8CA: sinewave <= 12'hD90;
        12'h8CB: sinewave <= 12'hD8D;
        12'h8CC: sinewave <= 12'hD8A;
        12'h8CD: sinewave <= 12'hD87;
        12'h8CE: sinewave <= 12'hD84;
        12'h8CF: sinewave <= 12'hD81;
        12'h8D0: sinewave <= 12'hD7E;
        12'h8D1: sinewave <= 12'hD7B;
        12'h8D2: sinewave <= 12'hD78;
        12'h8D3: sinewave <= 12'hD75;
        12'h8D4: sinewave <= 12'hD72;
        12'h8D5: sinewave <= 12'hD70;
        12'h8D6: sinewave <= 12'hD6D;
        12'h8D7: sinewave <= 12'hD6A;
        12'h8D8: sinewave <= 12'hD67;
        12'h8D9: sinewave <= 12'hD64;
        12'h8DA: sinewave <= 12'hD61;
        12'h8DB: sinewave <= 12'hD5E;
        12'h8DC: sinewave <= 12'hD5B;
        12'h8DD: sinewave <= 12'hD58;
        12'h8DE: sinewave <= 12'hD55;
        12'h8DF: sinewave <= 12'hD52;
        12'h8E0: sinewave <= 12'hD4F;
        12'h8E1: sinewave <= 12'hD4C;
        12'h8E2: sinewave <= 12'hD49;
        12'h8E3: sinewave <= 12'hD46;
        12'h8E4: sinewave <= 12'hD43;
        12'h8E5: sinewave <= 12'hD40;
        12'h8E6: sinewave <= 12'hD3D;
        12'h8E7: sinewave <= 12'hD3A;
        12'h8E8: sinewave <= 12'hD37;
        12'h8E9: sinewave <= 12'hD34;
        12'h8EA: sinewave <= 12'hD31;
        12'h8EB: sinewave <= 12'hD2E;
        12'h8EC: sinewave <= 12'hD2C;
        12'h8ED: sinewave <= 12'hD29;
        12'h8EE: sinewave <= 12'hD26;
        12'h8EF: sinewave <= 12'hD23;
        12'h8F0: sinewave <= 12'hD20;
        12'h8F1: sinewave <= 12'hD1D;
        12'h8F2: sinewave <= 12'hD1A;
        12'h8F3: sinewave <= 12'hD17;
        12'h8F4: sinewave <= 12'hD14;
        12'h8F5: sinewave <= 12'hD11;
        12'h8F6: sinewave <= 12'hD0E;
        12'h8F7: sinewave <= 12'hD0B;
        12'h8F8: sinewave <= 12'hD08;
        12'h8F9: sinewave <= 12'hD05;
        12'h8FA: sinewave <= 12'hD03;
        12'h8FB: sinewave <= 12'hD00;
        12'h8FC: sinewave <= 12'hCFD;
        12'h8FD: sinewave <= 12'hCFA;
        12'h8FE: sinewave <= 12'hCF7;
        12'h8FF: sinewave <= 12'hCF4;
        12'h900: sinewave <= 12'hCF1;
        12'h901: sinewave <= 12'hCEE;
        12'h902: sinewave <= 12'hCEB;
        12'h903: sinewave <= 12'hCE8;
        12'h904: sinewave <= 12'hCE6;
        12'h905: sinewave <= 12'hCE3;
        12'h906: sinewave <= 12'hCE0;
        12'h907: sinewave <= 12'hCDD;
        12'h908: sinewave <= 12'hCDA;
        12'h909: sinewave <= 12'hCD7;
        12'h90A: sinewave <= 12'hCD4;
        12'h90B: sinewave <= 12'hCD1;
        12'h90C: sinewave <= 12'hCCE;
        12'h90D: sinewave <= 12'hCCC;
        12'h90E: sinewave <= 12'hCC9;
        12'h90F: sinewave <= 12'hCC6;
        12'h910: sinewave <= 12'hCC3;
        12'h911: sinewave <= 12'hCC0;
        12'h912: sinewave <= 12'hCBD;
        12'h913: sinewave <= 12'hCBA;
        12'h914: sinewave <= 12'hCB8;
        12'h915: sinewave <= 12'hCB5;
        12'h916: sinewave <= 12'hCB2;
        12'h917: sinewave <= 12'hCAF;
        12'h918: sinewave <= 12'hCAC;
        12'h919: sinewave <= 12'hCA9;
        12'h91A: sinewave <= 12'hCA6;
        12'h91B: sinewave <= 12'hCA4;
        12'h91C: sinewave <= 12'hCA1;
        12'h91D: sinewave <= 12'hC9E;
        12'h91E: sinewave <= 12'hC9B;
        12'h91F: sinewave <= 12'hC98;
        12'h920: sinewave <= 12'hC95;
        12'h921: sinewave <= 12'hC92;
        12'h922: sinewave <= 12'hC90;
        12'h923: sinewave <= 12'hC8D;
        12'h924: sinewave <= 12'hC8A;
        12'h925: sinewave <= 12'hC87;
        12'h926: sinewave <= 12'hC84;
        12'h927: sinewave <= 12'hC81;
        12'h928: sinewave <= 12'hC7F;
        12'h929: sinewave <= 12'hC7C;
        12'h92A: sinewave <= 12'hC79;
        12'h92B: sinewave <= 12'hC76;
        12'h92C: sinewave <= 12'hC73;
        12'h92D: sinewave <= 12'hC71;
        12'h92E: sinewave <= 12'hC6E;
        12'h92F: sinewave <= 12'hC6B;
        12'h930: sinewave <= 12'hC68;
        12'h931: sinewave <= 12'hC65;
        12'h932: sinewave <= 12'hC63;
        12'h933: sinewave <= 12'hC60;
        12'h934: sinewave <= 12'hC5D;
        12'h935: sinewave <= 12'hC5A;
        12'h936: sinewave <= 12'hC57;
        12'h937: sinewave <= 12'hC55;
        12'h938: sinewave <= 12'hC52;
        12'h939: sinewave <= 12'hC4F;
        12'h93A: sinewave <= 12'hC4C;
        12'h93B: sinewave <= 12'hC49;
        12'h93C: sinewave <= 12'hC47;
        12'h93D: sinewave <= 12'hC44;
        12'h93E: sinewave <= 12'hC41;
        12'h93F: sinewave <= 12'hC3E;
        12'h940: sinewave <= 12'hC3C;
        12'h941: sinewave <= 12'hC39;
        12'h942: sinewave <= 12'hC36;
        12'h943: sinewave <= 12'hC33;
        12'h944: sinewave <= 12'hC30;
        12'h945: sinewave <= 12'hC2E;
        12'h946: sinewave <= 12'hC2B;
        12'h947: sinewave <= 12'hC28;
        12'h948: sinewave <= 12'hC25;
        12'h949: sinewave <= 12'hC23;
        12'h94A: sinewave <= 12'hC20;
        12'h94B: sinewave <= 12'hC1D;
        12'h94C: sinewave <= 12'hC1A;
        12'h94D: sinewave <= 12'hC18;
        12'h94E: sinewave <= 12'hC15;
        12'h94F: sinewave <= 12'hC12;
        12'h950: sinewave <= 12'hC10;
        12'h951: sinewave <= 12'hC0D;
        12'h952: sinewave <= 12'hC0A;
        12'h953: sinewave <= 12'hC07;
        12'h954: sinewave <= 12'hC05;
        12'h955: sinewave <= 12'hC02;
        12'h956: sinewave <= 12'hBFF;
        12'h957: sinewave <= 12'hBFC;
        12'h958: sinewave <= 12'hBFA;
        12'h959: sinewave <= 12'hBF7;
        12'h95A: sinewave <= 12'hBF4;
        12'h95B: sinewave <= 12'hBF2;
        12'h95C: sinewave <= 12'hBEF;
        12'h95D: sinewave <= 12'hBEC;
        12'h95E: sinewave <= 12'hBEA;
        12'h95F: sinewave <= 12'hBE7;
        12'h960: sinewave <= 12'hBE4;
        12'h961: sinewave <= 12'hBE1;
        12'h962: sinewave <= 12'hBDF;
        12'h963: sinewave <= 12'hBDC;
        12'h964: sinewave <= 12'hBD9;
        12'h965: sinewave <= 12'hBD7;
        12'h966: sinewave <= 12'hBD4;
        12'h967: sinewave <= 12'hBD1;
        12'h968: sinewave <= 12'hBCF;
        12'h969: sinewave <= 12'hBCC;
        12'h96A: sinewave <= 12'hBC9;
        12'h96B: sinewave <= 12'hBC7;
        12'h96C: sinewave <= 12'hBC4;
        12'h96D: sinewave <= 12'hBC1;
        12'h96E: sinewave <= 12'hBBF;
        12'h96F: sinewave <= 12'hBBC;
        12'h970: sinewave <= 12'hBB9;
        12'h971: sinewave <= 12'hBB7;
        12'h972: sinewave <= 12'hBB4;
        12'h973: sinewave <= 12'hBB1;
        12'h974: sinewave <= 12'hBAF;
        12'h975: sinewave <= 12'hBAC;
        12'h976: sinewave <= 12'hBA9;
        12'h977: sinewave <= 12'hBA7;
        12'h978: sinewave <= 12'hBA4;
        12'h979: sinewave <= 12'hBA2;
        12'h97A: sinewave <= 12'hB9F;
        12'h97B: sinewave <= 12'hB9C;
        12'h97C: sinewave <= 12'hB9A;
        12'h97D: sinewave <= 12'hB97;
        12'h97E: sinewave <= 12'hB94;
        12'h97F: sinewave <= 12'hB92;
        12'h980: sinewave <= 12'hB8F;
        12'h981: sinewave <= 12'hB8D;
        12'h982: sinewave <= 12'hB8A;
        12'h983: sinewave <= 12'hB87;
        12'h984: sinewave <= 12'hB85;
        12'h985: sinewave <= 12'hB82;
        12'h986: sinewave <= 12'hB80;
        12'h987: sinewave <= 12'hB7D;
        12'h988: sinewave <= 12'hB7A;
        12'h989: sinewave <= 12'hB78;
        12'h98A: sinewave <= 12'hB75;
        12'h98B: sinewave <= 12'hB73;
        12'h98C: sinewave <= 12'hB70;
        12'h98D: sinewave <= 12'hB6E;
        12'h98E: sinewave <= 12'hB6B;
        12'h98F: sinewave <= 12'hB68;
        12'h990: sinewave <= 12'hB66;
        12'h991: sinewave <= 12'hB63;
        12'h992: sinewave <= 12'hB61;
        12'h993: sinewave <= 12'hB5E;
        12'h994: sinewave <= 12'hB5C;
        12'h995: sinewave <= 12'hB59;
        12'h996: sinewave <= 12'hB56;
        12'h997: sinewave <= 12'hB54;
        12'h998: sinewave <= 12'hB51;
        12'h999: sinewave <= 12'hB4F;
        12'h99A: sinewave <= 12'hB4C;
        12'h99B: sinewave <= 12'hB4A;
        12'h99C: sinewave <= 12'hB47;
        12'h99D: sinewave <= 12'hB45;
        12'h99E: sinewave <= 12'hB42;
        12'h99F: sinewave <= 12'hB40;
        12'h9A0: sinewave <= 12'hB3D;
        12'h9A1: sinewave <= 12'hB3B;
        12'h9A2: sinewave <= 12'hB38;
        12'h9A3: sinewave <= 12'hB36;
        12'h9A4: sinewave <= 12'hB33;
        12'h9A5: sinewave <= 12'hB31;
        12'h9A6: sinewave <= 12'hB2E;
        12'h9A7: sinewave <= 12'hB2C;
        12'h9A8: sinewave <= 12'hB29;
        12'h9A9: sinewave <= 12'hB27;
        12'h9AA: sinewave <= 12'hB24;
        12'h9AB: sinewave <= 12'hB22;
        12'h9AC: sinewave <= 12'hB1F;
        12'h9AD: sinewave <= 12'hB1D;
        12'h9AE: sinewave <= 12'hB1A;
        12'h9AF: sinewave <= 12'hB18;
        12'h9B0: sinewave <= 12'hB15;
        12'h9B1: sinewave <= 12'hB13;
        12'h9B2: sinewave <= 12'hB10;
        12'h9B3: sinewave <= 12'hB0E;
        12'h9B4: sinewave <= 12'hB0B;
        12'h9B5: sinewave <= 12'hB09;
        12'h9B6: sinewave <= 12'hB06;
        12'h9B7: sinewave <= 12'hB04;
        12'h9B8: sinewave <= 12'hB01;
        12'h9B9: sinewave <= 12'hAFF;
        12'h9BA: sinewave <= 12'hAFD;
        12'h9BB: sinewave <= 12'hAFA;
        12'h9BC: sinewave <= 12'hAF8;
        12'h9BD: sinewave <= 12'hAF5;
        12'h9BE: sinewave <= 12'hAF3;
        12'h9BF: sinewave <= 12'hAF0;
        12'h9C0: sinewave <= 12'hAEE;
        12'h9C1: sinewave <= 12'hAEB;
        12'h9C2: sinewave <= 12'hAE9;
        12'h9C3: sinewave <= 12'hAE7;
        12'h9C4: sinewave <= 12'hAE4;
        12'h9C5: sinewave <= 12'hAE2;
        12'h9C6: sinewave <= 12'hADF;
        12'h9C7: sinewave <= 12'hADD;
        12'h9C8: sinewave <= 12'hADB;
        12'h9C9: sinewave <= 12'hAD8;
        12'h9CA: sinewave <= 12'hAD6;
        12'h9CB: sinewave <= 12'hAD3;
        12'h9CC: sinewave <= 12'hAD1;
        12'h9CD: sinewave <= 12'hACF;
        12'h9CE: sinewave <= 12'hACC;
        12'h9CF: sinewave <= 12'hACA;
        12'h9D0: sinewave <= 12'hAC7;
        12'h9D1: sinewave <= 12'hAC5;
        12'h9D2: sinewave <= 12'hAC3;
        12'h9D3: sinewave <= 12'hAC0;
        12'h9D4: sinewave <= 12'hABE;
        12'h9D5: sinewave <= 12'hABC;
        12'h9D6: sinewave <= 12'hAB9;
        12'h9D7: sinewave <= 12'hAB7;
        12'h9D8: sinewave <= 12'hAB5;
        12'h9D9: sinewave <= 12'hAB2;
        12'h9DA: sinewave <= 12'hAB0;
        12'h9DB: sinewave <= 12'hAAD;
        12'h9DC: sinewave <= 12'hAAB;
        12'h9DD: sinewave <= 12'hAA9;
        12'h9DE: sinewave <= 12'hAA6;
        12'h9DF: sinewave <= 12'hAA4;
        12'h9E0: sinewave <= 12'hAA2;
        12'h9E1: sinewave <= 12'hA9F;
        12'h9E2: sinewave <= 12'hA9D;
        12'h9E3: sinewave <= 12'hA9B;
        12'h9E4: sinewave <= 12'hA99;
        12'h9E5: sinewave <= 12'hA96;
        12'h9E6: sinewave <= 12'hA94;
        12'h9E7: sinewave <= 12'hA92;
        12'h9E8: sinewave <= 12'hA8F;
        12'h9E9: sinewave <= 12'hA8D;
        12'h9EA: sinewave <= 12'hA8B;
        12'h9EB: sinewave <= 12'hA88;
        12'h9EC: sinewave <= 12'hA86;
        12'h9ED: sinewave <= 12'hA84;
        12'h9EE: sinewave <= 12'hA82;
        12'h9EF: sinewave <= 12'hA7F;
        12'h9F0: sinewave <= 12'hA7D;
        12'h9F1: sinewave <= 12'hA7B;
        12'h9F2: sinewave <= 12'hA78;
        12'h9F3: sinewave <= 12'hA76;
        12'h9F4: sinewave <= 12'hA74;
        12'h9F5: sinewave <= 12'hA72;
        12'h9F6: sinewave <= 12'hA6F;
        12'h9F7: sinewave <= 12'hA6D;
        12'h9F8: sinewave <= 12'hA6B;
        12'h9F9: sinewave <= 12'hA69;
        12'h9FA: sinewave <= 12'hA66;
        12'h9FB: sinewave <= 12'hA64;
        12'h9FC: sinewave <= 12'hA62;
        12'h9FD: sinewave <= 12'hA60;
        12'h9FE: sinewave <= 12'hA5D;
        12'h9FF: sinewave <= 12'hA5B;
        12'hA00: sinewave <= 12'hA59;
        12'hA01: sinewave <= 12'hA57;
        12'hA02: sinewave <= 12'hA55;
        12'hA03: sinewave <= 12'hA52;
        12'hA04: sinewave <= 12'hA50;
        12'hA05: sinewave <= 12'hA4E;
        12'hA06: sinewave <= 12'hA4C;
        12'hA07: sinewave <= 12'hA4A;
        12'hA08: sinewave <= 12'hA47;
        12'hA09: sinewave <= 12'hA45;
        12'hA0A: sinewave <= 12'hA43;
        12'hA0B: sinewave <= 12'hA41;
        12'hA0C: sinewave <= 12'hA3F;
        12'hA0D: sinewave <= 12'hA3C;
        12'hA0E: sinewave <= 12'hA3A;
        12'hA0F: sinewave <= 12'hA38;
        12'hA10: sinewave <= 12'hA36;
        12'hA11: sinewave <= 12'hA34;
        12'hA12: sinewave <= 12'hA32;
        12'hA13: sinewave <= 12'hA2F;
        12'hA14: sinewave <= 12'hA2D;
        12'hA15: sinewave <= 12'hA2B;
        12'hA16: sinewave <= 12'hA29;
        12'hA17: sinewave <= 12'hA27;
        12'hA18: sinewave <= 12'hA25;
        12'hA19: sinewave <= 12'hA23;
        12'hA1A: sinewave <= 12'hA20;
        12'hA1B: sinewave <= 12'hA1E;
        12'hA1C: sinewave <= 12'hA1C;
        12'hA1D: sinewave <= 12'hA1A;
        12'hA1E: sinewave <= 12'hA18;
        12'hA1F: sinewave <= 12'hA16;
        12'hA20: sinewave <= 12'hA14;
        12'hA21: sinewave <= 12'hA12;
        12'hA22: sinewave <= 12'hA10;
        12'hA23: sinewave <= 12'hA0D;
        12'hA24: sinewave <= 12'hA0B;
        12'hA25: sinewave <= 12'hA09;
        12'hA26: sinewave <= 12'hA07;
        12'hA27: sinewave <= 12'hA05;
        12'hA28: sinewave <= 12'hA03;
        12'hA29: sinewave <= 12'hA01;
        12'hA2A: sinewave <= 12'h9FF;
        12'hA2B: sinewave <= 12'h9FD;
        12'hA2C: sinewave <= 12'h9FB;
        12'hA2D: sinewave <= 12'h9F9;
        12'hA2E: sinewave <= 12'h9F7;
        12'hA2F: sinewave <= 12'h9F5;
        12'hA30: sinewave <= 12'h9F2;
        12'hA31: sinewave <= 12'h9F0;
        12'hA32: sinewave <= 12'h9EE;
        12'hA33: sinewave <= 12'h9EC;
        12'hA34: sinewave <= 12'h9EA;
        12'hA35: sinewave <= 12'h9E8;
        12'hA36: sinewave <= 12'h9E6;
        12'hA37: sinewave <= 12'h9E4;
        12'hA38: sinewave <= 12'h9E2;
        12'hA39: sinewave <= 12'h9E0;
        12'hA3A: sinewave <= 12'h9DE;
        12'hA3B: sinewave <= 12'h9DC;
        12'hA3C: sinewave <= 12'h9DA;
        12'hA3D: sinewave <= 12'h9D8;
        12'hA3E: sinewave <= 12'h9D6;
        12'hA3F: sinewave <= 12'h9D4;
        12'hA40: sinewave <= 12'h9D2;
        12'hA41: sinewave <= 12'h9D0;
        12'hA42: sinewave <= 12'h9CE;
        12'hA43: sinewave <= 12'h9CC;
        12'hA44: sinewave <= 12'h9CA;
        12'hA45: sinewave <= 12'h9C8;
        12'hA46: sinewave <= 12'h9C6;
        12'hA47: sinewave <= 12'h9C4;
        12'hA48: sinewave <= 12'h9C2;
        12'hA49: sinewave <= 12'h9C0;
        12'hA4A: sinewave <= 12'h9BE;
        12'hA4B: sinewave <= 12'h9BC;
        12'hA4C: sinewave <= 12'h9BB;
        12'hA4D: sinewave <= 12'h9B9;
        12'hA4E: sinewave <= 12'h9B7;
        12'hA4F: sinewave <= 12'h9B5;
        12'hA50: sinewave <= 12'h9B3;
        12'hA51: sinewave <= 12'h9B1;
        12'hA52: sinewave <= 12'h9AF;
        12'hA53: sinewave <= 12'h9AD;
        12'hA54: sinewave <= 12'h9AB;
        12'hA55: sinewave <= 12'h9A9;
        12'hA56: sinewave <= 12'h9A7;
        12'hA57: sinewave <= 12'h9A5;
        12'hA58: sinewave <= 12'h9A3;
        12'hA59: sinewave <= 12'h9A2;
        12'hA5A: sinewave <= 12'h9A0;
        12'hA5B: sinewave <= 12'h99E;
        12'hA5C: sinewave <= 12'h99C;
        12'hA5D: sinewave <= 12'h99A;
        12'hA5E: sinewave <= 12'h998;
        12'hA5F: sinewave <= 12'h996;
        12'hA60: sinewave <= 12'h994;
        12'hA61: sinewave <= 12'h992;
        12'hA62: sinewave <= 12'h991;
        12'hA63: sinewave <= 12'h98F;
        12'hA64: sinewave <= 12'h98D;
        12'hA65: sinewave <= 12'h98B;
        12'hA66: sinewave <= 12'h989;
        12'hA67: sinewave <= 12'h987;
        12'hA68: sinewave <= 12'h985;
        12'hA69: sinewave <= 12'h984;
        12'hA6A: sinewave <= 12'h982;
        12'hA6B: sinewave <= 12'h980;
        12'hA6C: sinewave <= 12'h97E;
        12'hA6D: sinewave <= 12'h97C;
        12'hA6E: sinewave <= 12'h97B;
        12'hA6F: sinewave <= 12'h979;
        12'hA70: sinewave <= 12'h977;
        12'hA71: sinewave <= 12'h975;
        12'hA72: sinewave <= 12'h973;
        12'hA73: sinewave <= 12'h971;
        12'hA74: sinewave <= 12'h970;
        12'hA75: sinewave <= 12'h96E;
        12'hA76: sinewave <= 12'h96C;
        12'hA77: sinewave <= 12'h96A;
        12'hA78: sinewave <= 12'h969;
        12'hA79: sinewave <= 12'h967;
        12'hA7A: sinewave <= 12'h965;
        12'hA7B: sinewave <= 12'h963;
        12'hA7C: sinewave <= 12'h961;
        12'hA7D: sinewave <= 12'h960;
        12'hA7E: sinewave <= 12'h95E;
        12'hA7F: sinewave <= 12'h95C;
        12'hA80: sinewave <= 12'h95A;
        12'hA81: sinewave <= 12'h959;
        12'hA82: sinewave <= 12'h957;
        12'hA83: sinewave <= 12'h955;
        12'hA84: sinewave <= 12'h954;
        12'hA85: sinewave <= 12'h952;
        12'hA86: sinewave <= 12'h950;
        12'hA87: sinewave <= 12'h94E;
        12'hA88: sinewave <= 12'h94D;
        12'hA89: sinewave <= 12'h94B;
        12'hA8A: sinewave <= 12'h949;
        12'hA8B: sinewave <= 12'h948;
        12'hA8C: sinewave <= 12'h946;
        12'hA8D: sinewave <= 12'h944;
        12'hA8E: sinewave <= 12'h942;
        12'hA8F: sinewave <= 12'h941;
        12'hA90: sinewave <= 12'h93F;
        12'hA91: sinewave <= 12'h93D;
        12'hA92: sinewave <= 12'h93C;
        12'hA93: sinewave <= 12'h93A;
        12'hA94: sinewave <= 12'h938;
        12'hA95: sinewave <= 12'h937;
        12'hA96: sinewave <= 12'h935;
        12'hA97: sinewave <= 12'h933;
        12'hA98: sinewave <= 12'h932;
        12'hA99: sinewave <= 12'h930;
        12'hA9A: sinewave <= 12'h92E;
        12'hA9B: sinewave <= 12'h92D;
        12'hA9C: sinewave <= 12'h92B;
        12'hA9D: sinewave <= 12'h92A;
        12'hA9E: sinewave <= 12'h928;
        12'hA9F: sinewave <= 12'h926;
        12'hAA0: sinewave <= 12'h925;
        12'hAA1: sinewave <= 12'h923;
        12'hAA2: sinewave <= 12'h922;
        12'hAA3: sinewave <= 12'h920;
        12'hAA4: sinewave <= 12'h91E;
        12'hAA5: sinewave <= 12'h91D;
        12'hAA6: sinewave <= 12'h91B;
        12'hAA7: sinewave <= 12'h91A;
        12'hAA8: sinewave <= 12'h918;
        12'hAA9: sinewave <= 12'h916;
        12'hAAA: sinewave <= 12'h915;
        12'hAAB: sinewave <= 12'h913;
        12'hAAC: sinewave <= 12'h912;
        12'hAAD: sinewave <= 12'h910;
        12'hAAE: sinewave <= 12'h90F;
        12'hAAF: sinewave <= 12'h90D;
        12'hAB0: sinewave <= 12'h90B;
        12'hAB1: sinewave <= 12'h90A;
        12'hAB2: sinewave <= 12'h908;
        12'hAB3: sinewave <= 12'h907;
        12'hAB4: sinewave <= 12'h905;
        12'hAB5: sinewave <= 12'h904;
        12'hAB6: sinewave <= 12'h902;
        12'hAB7: sinewave <= 12'h901;
        12'hAB8: sinewave <= 12'h8FF;
        12'hAB9: sinewave <= 12'h8FE;
        12'hABA: sinewave <= 12'h8FC;
        12'hABB: sinewave <= 12'h8FB;
        12'hABC: sinewave <= 12'h8F9;
        12'hABD: sinewave <= 12'h8F8;
        12'hABE: sinewave <= 12'h8F6;
        12'hABF: sinewave <= 12'h8F5;
        12'hAC0: sinewave <= 12'h8F3;
        12'hAC1: sinewave <= 12'h8F2;
        12'hAC2: sinewave <= 12'h8F0;
        12'hAC3: sinewave <= 12'h8EF;
        12'hAC4: sinewave <= 12'h8ED;
        12'hAC5: sinewave <= 12'h8EC;
        12'hAC6: sinewave <= 12'h8EA;
        12'hAC7: sinewave <= 12'h8E9;
        12'hAC8: sinewave <= 12'h8E8;
        12'hAC9: sinewave <= 12'h8E6;
        12'hACA: sinewave <= 12'h8E5;
        12'hACB: sinewave <= 12'h8E3;
        12'hACC: sinewave <= 12'h8E2;
        12'hACD: sinewave <= 12'h8E0;
        12'hACE: sinewave <= 12'h8DF;
        12'hACF: sinewave <= 12'h8DD;
        12'hAD0: sinewave <= 12'h8DC;
        12'hAD1: sinewave <= 12'h8DB;
        12'hAD2: sinewave <= 12'h8D9;
        12'hAD3: sinewave <= 12'h8D8;
        12'hAD4: sinewave <= 12'h8D6;
        12'hAD5: sinewave <= 12'h8D5;
        12'hAD6: sinewave <= 12'h8D4;
        12'hAD7: sinewave <= 12'h8D2;
        12'hAD8: sinewave <= 12'h8D1;
        12'hAD9: sinewave <= 12'h8D0;
        12'hADA: sinewave <= 12'h8CE;
        12'hADB: sinewave <= 12'h8CD;
        12'hADC: sinewave <= 12'h8CB;
        12'hADD: sinewave <= 12'h8CA;
        12'hADE: sinewave <= 12'h8C9;
        12'hADF: sinewave <= 12'h8C7;
        12'hAE0: sinewave <= 12'h8C6;
        12'hAE1: sinewave <= 12'h8C5;
        12'hAE2: sinewave <= 12'h8C3;
        12'hAE3: sinewave <= 12'h8C2;
        12'hAE4: sinewave <= 12'h8C1;
        12'hAE5: sinewave <= 12'h8BF;
        12'hAE6: sinewave <= 12'h8BE;
        12'hAE7: sinewave <= 12'h8BD;
        12'hAE8: sinewave <= 12'h8BB;
        12'hAE9: sinewave <= 12'h8BA;
        12'hAEA: sinewave <= 12'h8B9;
        12'hAEB: sinewave <= 12'h8B8;
        12'hAEC: sinewave <= 12'h8B6;
        12'hAED: sinewave <= 12'h8B5;
        12'hAEE: sinewave <= 12'h8B4;
        12'hAEF: sinewave <= 12'h8B2;
        12'hAF0: sinewave <= 12'h8B1;
        12'hAF1: sinewave <= 12'h8B0;
        12'hAF2: sinewave <= 12'h8AF;
        12'hAF3: sinewave <= 12'h8AD;
        12'hAF4: sinewave <= 12'h8AC;
        12'hAF5: sinewave <= 12'h8AB;
        12'hAF6: sinewave <= 12'h8AA;
        12'hAF7: sinewave <= 12'h8A8;
        12'hAF8: sinewave <= 12'h8A7;
        12'hAF9: sinewave <= 12'h8A6;
        12'hAFA: sinewave <= 12'h8A5;
        12'hAFB: sinewave <= 12'h8A3;
        12'hAFC: sinewave <= 12'h8A2;
        12'hAFD: sinewave <= 12'h8A1;
        12'hAFE: sinewave <= 12'h8A0;
        12'hAFF: sinewave <= 12'h89F;
        12'hB00: sinewave <= 12'h89D;
        12'hB01: sinewave <= 12'h89C;
        12'hB02: sinewave <= 12'h89B;
        12'hB03: sinewave <= 12'h89A;
        12'hB04: sinewave <= 12'h899;
        12'hB05: sinewave <= 12'h897;
        12'hB06: sinewave <= 12'h896;
        12'hB07: sinewave <= 12'h895;
        12'hB08: sinewave <= 12'h894;
        12'hB09: sinewave <= 12'h893;
        12'hB0A: sinewave <= 12'h892;
        12'hB0B: sinewave <= 12'h890;
        12'hB0C: sinewave <= 12'h88F;
        12'hB0D: sinewave <= 12'h88E;
        12'hB0E: sinewave <= 12'h88D;
        12'hB0F: sinewave <= 12'h88C;
        12'hB10: sinewave <= 12'h88B;
        12'hB11: sinewave <= 12'h88A;
        12'hB12: sinewave <= 12'h888;
        12'hB13: sinewave <= 12'h887;
        12'hB14: sinewave <= 12'h886;
        12'hB15: sinewave <= 12'h885;
        12'hB16: sinewave <= 12'h884;
        12'hB17: sinewave <= 12'h883;
        12'hB18: sinewave <= 12'h882;
        12'hB19: sinewave <= 12'h881;
        12'hB1A: sinewave <= 12'h880;
        12'hB1B: sinewave <= 12'h87F;
        12'hB1C: sinewave <= 12'h87D;
        12'hB1D: sinewave <= 12'h87C;
        12'hB1E: sinewave <= 12'h87B;
        12'hB1F: sinewave <= 12'h87A;
        12'hB20: sinewave <= 12'h879;
        12'hB21: sinewave <= 12'h878;
        12'hB22: sinewave <= 12'h877;
        12'hB23: sinewave <= 12'h876;
        12'hB24: sinewave <= 12'h875;
        12'hB25: sinewave <= 12'h874;
        12'hB26: sinewave <= 12'h873;
        12'hB27: sinewave <= 12'h872;
        12'hB28: sinewave <= 12'h871;
        12'hB29: sinewave <= 12'h870;
        12'hB2A: sinewave <= 12'h86F;
        12'hB2B: sinewave <= 12'h86E;
        12'hB2C: sinewave <= 12'h86D;
        12'hB2D: sinewave <= 12'h86C;
        12'hB2E: sinewave <= 12'h86B;
        12'hB2F: sinewave <= 12'h86A;
        12'hB30: sinewave <= 12'h869;
        12'hB31: sinewave <= 12'h868;
        12'hB32: sinewave <= 12'h867;
        12'hB33: sinewave <= 12'h866;
        12'hB34: sinewave <= 12'h865;
        12'hB35: sinewave <= 12'h864;
        12'hB36: sinewave <= 12'h863;
        12'hB37: sinewave <= 12'h862;
        12'hB38: sinewave <= 12'h861;
        12'hB39: sinewave <= 12'h860;
        12'hB3A: sinewave <= 12'h85F;
        12'hB3B: sinewave <= 12'h85E;
        12'hB3C: sinewave <= 12'h85D;
        12'hB3D: sinewave <= 12'h85C;
        12'hB3E: sinewave <= 12'h85B;
        12'hB3F: sinewave <= 12'h85B;
        12'hB40: sinewave <= 12'h85A;
        12'hB41: sinewave <= 12'h859;
        12'hB42: sinewave <= 12'h858;
        12'hB43: sinewave <= 12'h857;
        12'hB44: sinewave <= 12'h856;
        12'hB45: sinewave <= 12'h855;
        12'hB46: sinewave <= 12'h854;
        12'hB47: sinewave <= 12'h853;
        12'hB48: sinewave <= 12'h852;
        12'hB49: sinewave <= 12'h852;
        12'hB4A: sinewave <= 12'h851;
        12'hB4B: sinewave <= 12'h850;
        12'hB4C: sinewave <= 12'h84F;
        12'hB4D: sinewave <= 12'h84E;
        12'hB4E: sinewave <= 12'h84D;
        12'hB4F: sinewave <= 12'h84C;
        12'hB50: sinewave <= 12'h84C;
        12'hB51: sinewave <= 12'h84B;
        12'hB52: sinewave <= 12'h84A;
        12'hB53: sinewave <= 12'h849;
        12'hB54: sinewave <= 12'h848;
        12'hB55: sinewave <= 12'h848;
        12'hB56: sinewave <= 12'h847;
        12'hB57: sinewave <= 12'h846;
        12'hB58: sinewave <= 12'h845;
        12'hB59: sinewave <= 12'h844;
        12'hB5A: sinewave <= 12'h844;
        12'hB5B: sinewave <= 12'h843;
        12'hB5C: sinewave <= 12'h842;
        12'hB5D: sinewave <= 12'h841;
        12'hB5E: sinewave <= 12'h840;
        12'hB5F: sinewave <= 12'h840;
        12'hB60: sinewave <= 12'h83F;
        12'hB61: sinewave <= 12'h83E;
        12'hB62: sinewave <= 12'h83D;
        12'hB63: sinewave <= 12'h83D;
        12'hB64: sinewave <= 12'h83C;
        12'hB65: sinewave <= 12'h83B;
        12'hB66: sinewave <= 12'h83A;
        12'hB67: sinewave <= 12'h83A;
        12'hB68: sinewave <= 12'h839;
        12'hB69: sinewave <= 12'h838;
        12'hB6A: sinewave <= 12'h837;
        12'hB6B: sinewave <= 12'h837;
        12'hB6C: sinewave <= 12'h836;
        12'hB6D: sinewave <= 12'h835;
        12'hB6E: sinewave <= 12'h835;
        12'hB6F: sinewave <= 12'h834;
        12'hB70: sinewave <= 12'h833;
        12'hB71: sinewave <= 12'h833;
        12'hB72: sinewave <= 12'h832;
        12'hB73: sinewave <= 12'h831;
        12'hB74: sinewave <= 12'h831;
        12'hB75: sinewave <= 12'h830;
        12'hB76: sinewave <= 12'h82F;
        12'hB77: sinewave <= 12'h82F;
        12'hB78: sinewave <= 12'h82E;
        12'hB79: sinewave <= 12'h82D;
        12'hB7A: sinewave <= 12'h82D;
        12'hB7B: sinewave <= 12'h82C;
        12'hB7C: sinewave <= 12'h82B;
        12'hB7D: sinewave <= 12'h82B;
        12'hB7E: sinewave <= 12'h82A;
        12'hB7F: sinewave <= 12'h829;
        12'hB80: sinewave <= 12'h829;
        12'hB81: sinewave <= 12'h828;
        12'hB82: sinewave <= 12'h828;
        12'hB83: sinewave <= 12'h827;
        12'hB84: sinewave <= 12'h826;
        12'hB85: sinewave <= 12'h826;
        12'hB86: sinewave <= 12'h825;
        12'hB87: sinewave <= 12'h825;
        12'hB88: sinewave <= 12'h824;
        12'hB89: sinewave <= 12'h824;
        12'hB8A: sinewave <= 12'h823;
        12'hB8B: sinewave <= 12'h822;
        12'hB8C: sinewave <= 12'h822;
        12'hB8D: sinewave <= 12'h821;
        12'hB8E: sinewave <= 12'h821;
        12'hB8F: sinewave <= 12'h820;
        12'hB90: sinewave <= 12'h820;
        12'hB91: sinewave <= 12'h81F;
        12'hB92: sinewave <= 12'h81F;
        12'hB93: sinewave <= 12'h81E;
        12'hB94: sinewave <= 12'h81E;
        12'hB95: sinewave <= 12'h81D;
        12'hB96: sinewave <= 12'h81D;
        12'hB97: sinewave <= 12'h81C;
        12'hB98: sinewave <= 12'h81B;
        12'hB99: sinewave <= 12'h81B;
        12'hB9A: sinewave <= 12'h81B;
        12'hB9B: sinewave <= 12'h81A;
        12'hB9C: sinewave <= 12'h81A;
        12'hB9D: sinewave <= 12'h819;
        12'hB9E: sinewave <= 12'h819;
        12'hB9F: sinewave <= 12'h818;
        12'hBA0: sinewave <= 12'h818;
        12'hBA1: sinewave <= 12'h817;
        12'hBA2: sinewave <= 12'h817;
        12'hBA3: sinewave <= 12'h816;
        12'hBA4: sinewave <= 12'h816;
        12'hBA5: sinewave <= 12'h815;
        12'hBA6: sinewave <= 12'h815;
        12'hBA7: sinewave <= 12'h815;
        12'hBA8: sinewave <= 12'h814;
        12'hBA9: sinewave <= 12'h814;
        12'hBAA: sinewave <= 12'h813;
        12'hBAB: sinewave <= 12'h813;
        12'hBAC: sinewave <= 12'h812;
        12'hBAD: sinewave <= 12'h812;
        12'hBAE: sinewave <= 12'h812;
        12'hBAF: sinewave <= 12'h811;
        12'hBB0: sinewave <= 12'h811;
        12'hBB1: sinewave <= 12'h811;
        12'hBB2: sinewave <= 12'h810;
        12'hBB3: sinewave <= 12'h810;
        12'hBB4: sinewave <= 12'h80F;
        12'hBB5: sinewave <= 12'h80F;
        12'hBB6: sinewave <= 12'h80F;
        12'hBB7: sinewave <= 12'h80E;
        12'hBB8: sinewave <= 12'h80E;
        12'hBB9: sinewave <= 12'h80E;
        12'hBBA: sinewave <= 12'h80D;
        12'hBBB: sinewave <= 12'h80D;
        12'hBBC: sinewave <= 12'h80D;
        12'hBBD: sinewave <= 12'h80C;
        12'hBBE: sinewave <= 12'h80C;
        12'hBBF: sinewave <= 12'h80C;
        12'hBC0: sinewave <= 12'h80B;
        12'hBC1: sinewave <= 12'h80B;
        12'hBC2: sinewave <= 12'h80B;
        12'hBC3: sinewave <= 12'h80A;
        12'hBC4: sinewave <= 12'h80A;
        12'hBC5: sinewave <= 12'h80A;
        12'hBC6: sinewave <= 12'h80A;
        12'hBC7: sinewave <= 12'h809;
        12'hBC8: sinewave <= 12'h809;
        12'hBC9: sinewave <= 12'h809;
        12'hBCA: sinewave <= 12'h809;
        12'hBCB: sinewave <= 12'h808;
        12'hBCC: sinewave <= 12'h808;
        12'hBCD: sinewave <= 12'h808;
        12'hBCE: sinewave <= 12'h808;
        12'hBCF: sinewave <= 12'h807;
        12'hBD0: sinewave <= 12'h807;
        12'hBD1: sinewave <= 12'h807;
        12'hBD2: sinewave <= 12'h807;
        12'hBD3: sinewave <= 12'h806;
        12'hBD4: sinewave <= 12'h806;
        12'hBD5: sinewave <= 12'h806;
        12'hBD6: sinewave <= 12'h806;
        12'hBD7: sinewave <= 12'h806;
        12'hBD8: sinewave <= 12'h805;
        12'hBD9: sinewave <= 12'h805;
        12'hBDA: sinewave <= 12'h805;
        12'hBDB: sinewave <= 12'h805;
        12'hBDC: sinewave <= 12'h805;
        12'hBDD: sinewave <= 12'h804;
        12'hBDE: sinewave <= 12'h804;
        12'hBDF: sinewave <= 12'h804;
        12'hBE0: sinewave <= 12'h804;
        12'hBE1: sinewave <= 12'h804;
        12'hBE2: sinewave <= 12'h804;
        12'hBE3: sinewave <= 12'h804;
        12'hBE4: sinewave <= 12'h803;
        12'hBE5: sinewave <= 12'h803;
        12'hBE6: sinewave <= 12'h803;
        12'hBE7: sinewave <= 12'h803;
        12'hBE8: sinewave <= 12'h803;
        12'hBE9: sinewave <= 12'h803;
        12'hBEA: sinewave <= 12'h803;
        12'hBEB: sinewave <= 12'h803;
        12'hBEC: sinewave <= 12'h802;
        12'hBED: sinewave <= 12'h802;
        12'hBEE: sinewave <= 12'h802;
        12'hBEF: sinewave <= 12'h802;
        12'hBF0: sinewave <= 12'h802;
        12'hBF1: sinewave <= 12'h802;
        12'hBF2: sinewave <= 12'h802;
        12'hBF3: sinewave <= 12'h802;
        12'hBF4: sinewave <= 12'h802;
        12'hBF5: sinewave <= 12'h802;
        12'hBF6: sinewave <= 12'h802;
        12'hBF7: sinewave <= 12'h802;
        12'hBF8: sinewave <= 12'h802;
        12'hBF9: sinewave <= 12'h802;
        12'hBFA: sinewave <= 12'h802;
        12'hBFB: sinewave <= 12'h802;
        12'hBFC: sinewave <= 12'h802;
        12'hBFD: sinewave <= 12'h802;
        12'hBFE: sinewave <= 12'h802;
        12'hBFF: sinewave <= 12'h802;
        12'hC00: sinewave <= 12'h801;
        12'hC01: sinewave <= 12'h802;
        12'hC02: sinewave <= 12'h802;
        12'hC03: sinewave <= 12'h802;
        12'hC04: sinewave <= 12'h802;
        12'hC05: sinewave <= 12'h802;
        12'hC06: sinewave <= 12'h802;
        12'hC07: sinewave <= 12'h802;
        12'hC08: sinewave <= 12'h802;
        12'hC09: sinewave <= 12'h802;
        12'hC0A: sinewave <= 12'h802;
        12'hC0B: sinewave <= 12'h802;
        12'hC0C: sinewave <= 12'h802;
        12'hC0D: sinewave <= 12'h802;
        12'hC0E: sinewave <= 12'h802;
        12'hC0F: sinewave <= 12'h802;
        12'hC10: sinewave <= 12'h802;
        12'hC11: sinewave <= 12'h802;
        12'hC12: sinewave <= 12'h802;
        12'hC13: sinewave <= 12'h802;
        12'hC14: sinewave <= 12'h802;
        12'hC15: sinewave <= 12'h803;
        12'hC16: sinewave <= 12'h803;
        12'hC17: sinewave <= 12'h803;
        12'hC18: sinewave <= 12'h803;
        12'hC19: sinewave <= 12'h803;
        12'hC1A: sinewave <= 12'h803;
        12'hC1B: sinewave <= 12'h803;
        12'hC1C: sinewave <= 12'h803;
        12'hC1D: sinewave <= 12'h804;
        12'hC1E: sinewave <= 12'h804;
        12'hC1F: sinewave <= 12'h804;
        12'hC20: sinewave <= 12'h804;
        12'hC21: sinewave <= 12'h804;
        12'hC22: sinewave <= 12'h804;
        12'hC23: sinewave <= 12'h804;
        12'hC24: sinewave <= 12'h805;
        12'hC25: sinewave <= 12'h805;
        12'hC26: sinewave <= 12'h805;
        12'hC27: sinewave <= 12'h805;
        12'hC28: sinewave <= 12'h805;
        12'hC29: sinewave <= 12'h806;
        12'hC2A: sinewave <= 12'h806;
        12'hC2B: sinewave <= 12'h806;
        12'hC2C: sinewave <= 12'h806;
        12'hC2D: sinewave <= 12'h806;
        12'hC2E: sinewave <= 12'h807;
        12'hC2F: sinewave <= 12'h807;
        12'hC30: sinewave <= 12'h807;
        12'hC31: sinewave <= 12'h807;
        12'hC32: sinewave <= 12'h808;
        12'hC33: sinewave <= 12'h808;
        12'hC34: sinewave <= 12'h808;
        12'hC35: sinewave <= 12'h808;
        12'hC36: sinewave <= 12'h809;
        12'hC37: sinewave <= 12'h809;
        12'hC38: sinewave <= 12'h809;
        12'hC39: sinewave <= 12'h809;
        12'hC3A: sinewave <= 12'h80A;
        12'hC3B: sinewave <= 12'h80A;
        12'hC3C: sinewave <= 12'h80A;
        12'hC3D: sinewave <= 12'h80A;
        12'hC3E: sinewave <= 12'h80B;
        12'hC3F: sinewave <= 12'h80B;
        12'hC40: sinewave <= 12'h80B;
        12'hC41: sinewave <= 12'h80C;
        12'hC42: sinewave <= 12'h80C;
        12'hC43: sinewave <= 12'h80C;
        12'hC44: sinewave <= 12'h80D;
        12'hC45: sinewave <= 12'h80D;
        12'hC46: sinewave <= 12'h80D;
        12'hC47: sinewave <= 12'h80E;
        12'hC48: sinewave <= 12'h80E;
        12'hC49: sinewave <= 12'h80E;
        12'hC4A: sinewave <= 12'h80F;
        12'hC4B: sinewave <= 12'h80F;
        12'hC4C: sinewave <= 12'h80F;
        12'hC4D: sinewave <= 12'h810;
        12'hC4E: sinewave <= 12'h810;
        12'hC4F: sinewave <= 12'h811;
        12'hC50: sinewave <= 12'h811;
        12'hC51: sinewave <= 12'h811;
        12'hC52: sinewave <= 12'h812;
        12'hC53: sinewave <= 12'h812;
        12'hC54: sinewave <= 12'h812;
        12'hC55: sinewave <= 12'h813;
        12'hC56: sinewave <= 12'h813;
        12'hC57: sinewave <= 12'h814;
        12'hC58: sinewave <= 12'h814;
        12'hC59: sinewave <= 12'h815;
        12'hC5A: sinewave <= 12'h815;
        12'hC5B: sinewave <= 12'h815;
        12'hC5C: sinewave <= 12'h816;
        12'hC5D: sinewave <= 12'h816;
        12'hC5E: sinewave <= 12'h817;
        12'hC5F: sinewave <= 12'h817;
        12'hC60: sinewave <= 12'h818;
        12'hC61: sinewave <= 12'h818;
        12'hC62: sinewave <= 12'h819;
        12'hC63: sinewave <= 12'h819;
        12'hC64: sinewave <= 12'h81A;
        12'hC65: sinewave <= 12'h81A;
        12'hC66: sinewave <= 12'h81B;
        12'hC67: sinewave <= 12'h81B;
        12'hC68: sinewave <= 12'h81B;
        12'hC69: sinewave <= 12'h81C;
        12'hC6A: sinewave <= 12'h81D;
        12'hC6B: sinewave <= 12'h81D;
        12'hC6C: sinewave <= 12'h81E;
        12'hC6D: sinewave <= 12'h81E;
        12'hC6E: sinewave <= 12'h81F;
        12'hC6F: sinewave <= 12'h81F;
        12'hC70: sinewave <= 12'h820;
        12'hC71: sinewave <= 12'h820;
        12'hC72: sinewave <= 12'h821;
        12'hC73: sinewave <= 12'h821;
        12'hC74: sinewave <= 12'h822;
        12'hC75: sinewave <= 12'h822;
        12'hC76: sinewave <= 12'h823;
        12'hC77: sinewave <= 12'h824;
        12'hC78: sinewave <= 12'h824;
        12'hC79: sinewave <= 12'h825;
        12'hC7A: sinewave <= 12'h825;
        12'hC7B: sinewave <= 12'h826;
        12'hC7C: sinewave <= 12'h826;
        12'hC7D: sinewave <= 12'h827;
        12'hC7E: sinewave <= 12'h828;
        12'hC7F: sinewave <= 12'h828;
        12'hC80: sinewave <= 12'h829;
        12'hC81: sinewave <= 12'h829;
        12'hC82: sinewave <= 12'h82A;
        12'hC83: sinewave <= 12'h82B;
        12'hC84: sinewave <= 12'h82B;
        12'hC85: sinewave <= 12'h82C;
        12'hC86: sinewave <= 12'h82D;
        12'hC87: sinewave <= 12'h82D;
        12'hC88: sinewave <= 12'h82E;
        12'hC89: sinewave <= 12'h82F;
        12'hC8A: sinewave <= 12'h82F;
        12'hC8B: sinewave <= 12'h830;
        12'hC8C: sinewave <= 12'h831;
        12'hC8D: sinewave <= 12'h831;
        12'hC8E: sinewave <= 12'h832;
        12'hC8F: sinewave <= 12'h833;
        12'hC90: sinewave <= 12'h833;
        12'hC91: sinewave <= 12'h834;
        12'hC92: sinewave <= 12'h835;
        12'hC93: sinewave <= 12'h835;
        12'hC94: sinewave <= 12'h836;
        12'hC95: sinewave <= 12'h837;
        12'hC96: sinewave <= 12'h837;
        12'hC97: sinewave <= 12'h838;
        12'hC98: sinewave <= 12'h839;
        12'hC99: sinewave <= 12'h83A;
        12'hC9A: sinewave <= 12'h83A;
        12'hC9B: sinewave <= 12'h83B;
        12'hC9C: sinewave <= 12'h83C;
        12'hC9D: sinewave <= 12'h83D;
        12'hC9E: sinewave <= 12'h83D;
        12'hC9F: sinewave <= 12'h83E;
        12'hCA0: sinewave <= 12'h83F;
        12'hCA1: sinewave <= 12'h840;
        12'hCA2: sinewave <= 12'h840;
        12'hCA3: sinewave <= 12'h841;
        12'hCA4: sinewave <= 12'h842;
        12'hCA5: sinewave <= 12'h843;
        12'hCA6: sinewave <= 12'h844;
        12'hCA7: sinewave <= 12'h844;
        12'hCA8: sinewave <= 12'h845;
        12'hCA9: sinewave <= 12'h846;
        12'hCAA: sinewave <= 12'h847;
        12'hCAB: sinewave <= 12'h848;
        12'hCAC: sinewave <= 12'h848;
        12'hCAD: sinewave <= 12'h849;
        12'hCAE: sinewave <= 12'h84A;
        12'hCAF: sinewave <= 12'h84B;
        12'hCB0: sinewave <= 12'h84C;
        12'hCB1: sinewave <= 12'h84C;
        12'hCB2: sinewave <= 12'h84D;
        12'hCB3: sinewave <= 12'h84E;
        12'hCB4: sinewave <= 12'h84F;
        12'hCB5: sinewave <= 12'h850;
        12'hCB6: sinewave <= 12'h851;
        12'hCB7: sinewave <= 12'h852;
        12'hCB8: sinewave <= 12'h852;
        12'hCB9: sinewave <= 12'h853;
        12'hCBA: sinewave <= 12'h854;
        12'hCBB: sinewave <= 12'h855;
        12'hCBC: sinewave <= 12'h856;
        12'hCBD: sinewave <= 12'h857;
        12'hCBE: sinewave <= 12'h858;
        12'hCBF: sinewave <= 12'h859;
        12'hCC0: sinewave <= 12'h85A;
        12'hCC1: sinewave <= 12'h85B;
        12'hCC2: sinewave <= 12'h85B;
        12'hCC3: sinewave <= 12'h85C;
        12'hCC4: sinewave <= 12'h85D;
        12'hCC5: sinewave <= 12'h85E;
        12'hCC6: sinewave <= 12'h85F;
        12'hCC7: sinewave <= 12'h860;
        12'hCC8: sinewave <= 12'h861;
        12'hCC9: sinewave <= 12'h862;
        12'hCCA: sinewave <= 12'h863;
        12'hCCB: sinewave <= 12'h864;
        12'hCCC: sinewave <= 12'h865;
        12'hCCD: sinewave <= 12'h866;
        12'hCCE: sinewave <= 12'h867;
        12'hCCF: sinewave <= 12'h868;
        12'hCD0: sinewave <= 12'h869;
        12'hCD1: sinewave <= 12'h86A;
        12'hCD2: sinewave <= 12'h86B;
        12'hCD3: sinewave <= 12'h86C;
        12'hCD4: sinewave <= 12'h86D;
        12'hCD5: sinewave <= 12'h86E;
        12'hCD6: sinewave <= 12'h86F;
        12'hCD7: sinewave <= 12'h870;
        12'hCD8: sinewave <= 12'h871;
        12'hCD9: sinewave <= 12'h872;
        12'hCDA: sinewave <= 12'h873;
        12'hCDB: sinewave <= 12'h874;
        12'hCDC: sinewave <= 12'h875;
        12'hCDD: sinewave <= 12'h876;
        12'hCDE: sinewave <= 12'h877;
        12'hCDF: sinewave <= 12'h878;
        12'hCE0: sinewave <= 12'h879;
        12'hCE1: sinewave <= 12'h87A;
        12'hCE2: sinewave <= 12'h87B;
        12'hCE3: sinewave <= 12'h87C;
        12'hCE4: sinewave <= 12'h87D;
        12'hCE5: sinewave <= 12'h87F;
        12'hCE6: sinewave <= 12'h880;
        12'hCE7: sinewave <= 12'h881;
        12'hCE8: sinewave <= 12'h882;
        12'hCE9: sinewave <= 12'h883;
        12'hCEA: sinewave <= 12'h884;
        12'hCEB: sinewave <= 12'h885;
        12'hCEC: sinewave <= 12'h886;
        12'hCED: sinewave <= 12'h887;
        12'hCEE: sinewave <= 12'h888;
        12'hCEF: sinewave <= 12'h88A;
        12'hCF0: sinewave <= 12'h88B;
        12'hCF1: sinewave <= 12'h88C;
        12'hCF2: sinewave <= 12'h88D;
        12'hCF3: sinewave <= 12'h88E;
        12'hCF4: sinewave <= 12'h88F;
        12'hCF5: sinewave <= 12'h890;
        12'hCF6: sinewave <= 12'h892;
        12'hCF7: sinewave <= 12'h893;
        12'hCF8: sinewave <= 12'h894;
        12'hCF9: sinewave <= 12'h895;
        12'hCFA: sinewave <= 12'h896;
        12'hCFB: sinewave <= 12'h897;
        12'hCFC: sinewave <= 12'h899;
        12'hCFD: sinewave <= 12'h89A;
        12'hCFE: sinewave <= 12'h89B;
        12'hCFF: sinewave <= 12'h89C;
        12'hD00: sinewave <= 12'h89D;
        12'hD01: sinewave <= 12'h89F;
        12'hD02: sinewave <= 12'h8A0;
        12'hD03: sinewave <= 12'h8A1;
        12'hD04: sinewave <= 12'h8A2;
        12'hD05: sinewave <= 12'h8A3;
        12'hD06: sinewave <= 12'h8A5;
        12'hD07: sinewave <= 12'h8A6;
        12'hD08: sinewave <= 12'h8A7;
        12'hD09: sinewave <= 12'h8A8;
        12'hD0A: sinewave <= 12'h8AA;
        12'hD0B: sinewave <= 12'h8AB;
        12'hD0C: sinewave <= 12'h8AC;
        12'hD0D: sinewave <= 12'h8AD;
        12'hD0E: sinewave <= 12'h8AF;
        12'hD0F: sinewave <= 12'h8B0;
        12'hD10: sinewave <= 12'h8B1;
        12'hD11: sinewave <= 12'h8B2;
        12'hD12: sinewave <= 12'h8B4;
        12'hD13: sinewave <= 12'h8B5;
        12'hD14: sinewave <= 12'h8B6;
        12'hD15: sinewave <= 12'h8B8;
        12'hD16: sinewave <= 12'h8B9;
        12'hD17: sinewave <= 12'h8BA;
        12'hD18: sinewave <= 12'h8BB;
        12'hD19: sinewave <= 12'h8BD;
        12'hD1A: sinewave <= 12'h8BE;
        12'hD1B: sinewave <= 12'h8BF;
        12'hD1C: sinewave <= 12'h8C1;
        12'hD1D: sinewave <= 12'h8C2;
        12'hD1E: sinewave <= 12'h8C3;
        12'hD1F: sinewave <= 12'h8C5;
        12'hD20: sinewave <= 12'h8C6;
        12'hD21: sinewave <= 12'h8C7;
        12'hD22: sinewave <= 12'h8C9;
        12'hD23: sinewave <= 12'h8CA;
        12'hD24: sinewave <= 12'h8CB;
        12'hD25: sinewave <= 12'h8CD;
        12'hD26: sinewave <= 12'h8CE;
        12'hD27: sinewave <= 12'h8D0;
        12'hD28: sinewave <= 12'h8D1;
        12'hD29: sinewave <= 12'h8D2;
        12'hD2A: sinewave <= 12'h8D4;
        12'hD2B: sinewave <= 12'h8D5;
        12'hD2C: sinewave <= 12'h8D6;
        12'hD2D: sinewave <= 12'h8D8;
        12'hD2E: sinewave <= 12'h8D9;
        12'hD2F: sinewave <= 12'h8DB;
        12'hD30: sinewave <= 12'h8DC;
        12'hD31: sinewave <= 12'h8DD;
        12'hD32: sinewave <= 12'h8DF;
        12'hD33: sinewave <= 12'h8E0;
        12'hD34: sinewave <= 12'h8E2;
        12'hD35: sinewave <= 12'h8E3;
        12'hD36: sinewave <= 12'h8E5;
        12'hD37: sinewave <= 12'h8E6;
        12'hD38: sinewave <= 12'h8E8;
        12'hD39: sinewave <= 12'h8E9;
        12'hD3A: sinewave <= 12'h8EA;
        12'hD3B: sinewave <= 12'h8EC;
        12'hD3C: sinewave <= 12'h8ED;
        12'hD3D: sinewave <= 12'h8EF;
        12'hD3E: sinewave <= 12'h8F0;
        12'hD3F: sinewave <= 12'h8F2;
        12'hD40: sinewave <= 12'h8F3;
        12'hD41: sinewave <= 12'h8F5;
        12'hD42: sinewave <= 12'h8F6;
        12'hD43: sinewave <= 12'h8F8;
        12'hD44: sinewave <= 12'h8F9;
        12'hD45: sinewave <= 12'h8FB;
        12'hD46: sinewave <= 12'h8FC;
        12'hD47: sinewave <= 12'h8FE;
        12'hD48: sinewave <= 12'h8FF;
        12'hD49: sinewave <= 12'h901;
        12'hD4A: sinewave <= 12'h902;
        12'hD4B: sinewave <= 12'h904;
        12'hD4C: sinewave <= 12'h905;
        12'hD4D: sinewave <= 12'h907;
        12'hD4E: sinewave <= 12'h908;
        12'hD4F: sinewave <= 12'h90A;
        12'hD50: sinewave <= 12'h90B;
        12'hD51: sinewave <= 12'h90D;
        12'hD52: sinewave <= 12'h90F;
        12'hD53: sinewave <= 12'h910;
        12'hD54: sinewave <= 12'h912;
        12'hD55: sinewave <= 12'h913;
        12'hD56: sinewave <= 12'h915;
        12'hD57: sinewave <= 12'h916;
        12'hD58: sinewave <= 12'h918;
        12'hD59: sinewave <= 12'h91A;
        12'hD5A: sinewave <= 12'h91B;
        12'hD5B: sinewave <= 12'h91D;
        12'hD5C: sinewave <= 12'h91E;
        12'hD5D: sinewave <= 12'h920;
        12'hD5E: sinewave <= 12'h922;
        12'hD5F: sinewave <= 12'h923;
        12'hD60: sinewave <= 12'h925;
        12'hD61: sinewave <= 12'h926;
        12'hD62: sinewave <= 12'h928;
        12'hD63: sinewave <= 12'h92A;
        12'hD64: sinewave <= 12'h92B;
        12'hD65: sinewave <= 12'h92D;
        12'hD66: sinewave <= 12'h92E;
        12'hD67: sinewave <= 12'h930;
        12'hD68: sinewave <= 12'h932;
        12'hD69: sinewave <= 12'h933;
        12'hD6A: sinewave <= 12'h935;
        12'hD6B: sinewave <= 12'h937;
        12'hD6C: sinewave <= 12'h938;
        12'hD6D: sinewave <= 12'h93A;
        12'hD6E: sinewave <= 12'h93C;
        12'hD6F: sinewave <= 12'h93D;
        12'hD70: sinewave <= 12'h93F;
        12'hD71: sinewave <= 12'h941;
        12'hD72: sinewave <= 12'h942;
        12'hD73: sinewave <= 12'h944;
        12'hD74: sinewave <= 12'h946;
        12'hD75: sinewave <= 12'h948;
        12'hD76: sinewave <= 12'h949;
        12'hD77: sinewave <= 12'h94B;
        12'hD78: sinewave <= 12'h94D;
        12'hD79: sinewave <= 12'h94E;
        12'hD7A: sinewave <= 12'h950;
        12'hD7B: sinewave <= 12'h952;
        12'hD7C: sinewave <= 12'h954;
        12'hD7D: sinewave <= 12'h955;
        12'hD7E: sinewave <= 12'h957;
        12'hD7F: sinewave <= 12'h959;
        12'hD80: sinewave <= 12'h95A;
        12'hD81: sinewave <= 12'h95C;
        12'hD82: sinewave <= 12'h95E;
        12'hD83: sinewave <= 12'h960;
        12'hD84: sinewave <= 12'h961;
        12'hD85: sinewave <= 12'h963;
        12'hD86: sinewave <= 12'h965;
        12'hD87: sinewave <= 12'h967;
        12'hD88: sinewave <= 12'h969;
        12'hD89: sinewave <= 12'h96A;
        12'hD8A: sinewave <= 12'h96C;
        12'hD8B: sinewave <= 12'h96E;
        12'hD8C: sinewave <= 12'h970;
        12'hD8D: sinewave <= 12'h971;
        12'hD8E: sinewave <= 12'h973;
        12'hD8F: sinewave <= 12'h975;
        12'hD90: sinewave <= 12'h977;
        12'hD91: sinewave <= 12'h979;
        12'hD92: sinewave <= 12'h97B;
        12'hD93: sinewave <= 12'h97C;
        12'hD94: sinewave <= 12'h97E;
        12'hD95: sinewave <= 12'h980;
        12'hD96: sinewave <= 12'h982;
        12'hD97: sinewave <= 12'h984;
        12'hD98: sinewave <= 12'h985;
        12'hD99: sinewave <= 12'h987;
        12'hD9A: sinewave <= 12'h989;
        12'hD9B: sinewave <= 12'h98B;
        12'hD9C: sinewave <= 12'h98D;
        12'hD9D: sinewave <= 12'h98F;
        12'hD9E: sinewave <= 12'h991;
        12'hD9F: sinewave <= 12'h992;
        12'hDA0: sinewave <= 12'h994;
        12'hDA1: sinewave <= 12'h996;
        12'hDA2: sinewave <= 12'h998;
        12'hDA3: sinewave <= 12'h99A;
        12'hDA4: sinewave <= 12'h99C;
        12'hDA5: sinewave <= 12'h99E;
        12'hDA6: sinewave <= 12'h9A0;
        12'hDA7: sinewave <= 12'h9A2;
        12'hDA8: sinewave <= 12'h9A3;
        12'hDA9: sinewave <= 12'h9A5;
        12'hDAA: sinewave <= 12'h9A7;
        12'hDAB: sinewave <= 12'h9A9;
        12'hDAC: sinewave <= 12'h9AB;
        12'hDAD: sinewave <= 12'h9AD;
        12'hDAE: sinewave <= 12'h9AF;
        12'hDAF: sinewave <= 12'h9B1;
        12'hDB0: sinewave <= 12'h9B3;
        12'hDB1: sinewave <= 12'h9B5;
        12'hDB2: sinewave <= 12'h9B7;
        12'hDB3: sinewave <= 12'h9B9;
        12'hDB4: sinewave <= 12'h9BB;
        12'hDB5: sinewave <= 12'h9BC;
        12'hDB6: sinewave <= 12'h9BE;
        12'hDB7: sinewave <= 12'h9C0;
        12'hDB8: sinewave <= 12'h9C2;
        12'hDB9: sinewave <= 12'h9C4;
        12'hDBA: sinewave <= 12'h9C6;
        12'hDBB: sinewave <= 12'h9C8;
        12'hDBC: sinewave <= 12'h9CA;
        12'hDBD: sinewave <= 12'h9CC;
        12'hDBE: sinewave <= 12'h9CE;
        12'hDBF: sinewave <= 12'h9D0;
        12'hDC0: sinewave <= 12'h9D2;
        12'hDC1: sinewave <= 12'h9D4;
        12'hDC2: sinewave <= 12'h9D6;
        12'hDC3: sinewave <= 12'h9D8;
        12'hDC4: sinewave <= 12'h9DA;
        12'hDC5: sinewave <= 12'h9DC;
        12'hDC6: sinewave <= 12'h9DE;
        12'hDC7: sinewave <= 12'h9E0;
        12'hDC8: sinewave <= 12'h9E2;
        12'hDC9: sinewave <= 12'h9E4;
        12'hDCA: sinewave <= 12'h9E6;
        12'hDCB: sinewave <= 12'h9E8;
        12'hDCC: sinewave <= 12'h9EA;
        12'hDCD: sinewave <= 12'h9EC;
        12'hDCE: sinewave <= 12'h9EE;
        12'hDCF: sinewave <= 12'h9F0;
        12'hDD0: sinewave <= 12'h9F2;
        12'hDD1: sinewave <= 12'h9F5;
        12'hDD2: sinewave <= 12'h9F7;
        12'hDD3: sinewave <= 12'h9F9;
        12'hDD4: sinewave <= 12'h9FB;
        12'hDD5: sinewave <= 12'h9FD;
        12'hDD6: sinewave <= 12'h9FF;
        12'hDD7: sinewave <= 12'hA01;
        12'hDD8: sinewave <= 12'hA03;
        12'hDD9: sinewave <= 12'hA05;
        12'hDDA: sinewave <= 12'hA07;
        12'hDDB: sinewave <= 12'hA09;
        12'hDDC: sinewave <= 12'hA0B;
        12'hDDD: sinewave <= 12'hA0D;
        12'hDDE: sinewave <= 12'hA10;
        12'hDDF: sinewave <= 12'hA12;
        12'hDE0: sinewave <= 12'hA14;
        12'hDE1: sinewave <= 12'hA16;
        12'hDE2: sinewave <= 12'hA18;
        12'hDE3: sinewave <= 12'hA1A;
        12'hDE4: sinewave <= 12'hA1C;
        12'hDE5: sinewave <= 12'hA1E;
        12'hDE6: sinewave <= 12'hA20;
        12'hDE7: sinewave <= 12'hA23;
        12'hDE8: sinewave <= 12'hA25;
        12'hDE9: sinewave <= 12'hA27;
        12'hDEA: sinewave <= 12'hA29;
        12'hDEB: sinewave <= 12'hA2B;
        12'hDEC: sinewave <= 12'hA2D;
        12'hDED: sinewave <= 12'hA2F;
        12'hDEE: sinewave <= 12'hA32;
        12'hDEF: sinewave <= 12'hA34;
        12'hDF0: sinewave <= 12'hA36;
        12'hDF1: sinewave <= 12'hA38;
        12'hDF2: sinewave <= 12'hA3A;
        12'hDF3: sinewave <= 12'hA3C;
        12'hDF4: sinewave <= 12'hA3F;
        12'hDF5: sinewave <= 12'hA41;
        12'hDF6: sinewave <= 12'hA43;
        12'hDF7: sinewave <= 12'hA45;
        12'hDF8: sinewave <= 12'hA47;
        12'hDF9: sinewave <= 12'hA4A;
        12'hDFA: sinewave <= 12'hA4C;
        12'hDFB: sinewave <= 12'hA4E;
        12'hDFC: sinewave <= 12'hA50;
        12'hDFD: sinewave <= 12'hA52;
        12'hDFE: sinewave <= 12'hA55;
        12'hDFF: sinewave <= 12'hA57;
        12'hE00: sinewave <= 12'hA59;
        12'hE01: sinewave <= 12'hA5B;
        12'hE02: sinewave <= 12'hA5D;
        12'hE03: sinewave <= 12'hA60;
        12'hE04: sinewave <= 12'hA62;
        12'hE05: sinewave <= 12'hA64;
        12'hE06: sinewave <= 12'hA66;
        12'hE07: sinewave <= 12'hA69;
        12'hE08: sinewave <= 12'hA6B;
        12'hE09: sinewave <= 12'hA6D;
        12'hE0A: sinewave <= 12'hA6F;
        12'hE0B: sinewave <= 12'hA72;
        12'hE0C: sinewave <= 12'hA74;
        12'hE0D: sinewave <= 12'hA76;
        12'hE0E: sinewave <= 12'hA78;
        12'hE0F: sinewave <= 12'hA7B;
        12'hE10: sinewave <= 12'hA7D;
        12'hE11: sinewave <= 12'hA7F;
        12'hE12: sinewave <= 12'hA82;
        12'hE13: sinewave <= 12'hA84;
        12'hE14: sinewave <= 12'hA86;
        12'hE15: sinewave <= 12'hA88;
        12'hE16: sinewave <= 12'hA8B;
        12'hE17: sinewave <= 12'hA8D;
        12'hE18: sinewave <= 12'hA8F;
        12'hE19: sinewave <= 12'hA92;
        12'hE1A: sinewave <= 12'hA94;
        12'hE1B: sinewave <= 12'hA96;
        12'hE1C: sinewave <= 12'hA99;
        12'hE1D: sinewave <= 12'hA9B;
        12'hE1E: sinewave <= 12'hA9D;
        12'hE1F: sinewave <= 12'hA9F;
        12'hE20: sinewave <= 12'hAA2;
        12'hE21: sinewave <= 12'hAA4;
        12'hE22: sinewave <= 12'hAA6;
        12'hE23: sinewave <= 12'hAA9;
        12'hE24: sinewave <= 12'hAAB;
        12'hE25: sinewave <= 12'hAAD;
        12'hE26: sinewave <= 12'hAB0;
        12'hE27: sinewave <= 12'hAB2;
        12'hE28: sinewave <= 12'hAB5;
        12'hE29: sinewave <= 12'hAB7;
        12'hE2A: sinewave <= 12'hAB9;
        12'hE2B: sinewave <= 12'hABC;
        12'hE2C: sinewave <= 12'hABE;
        12'hE2D: sinewave <= 12'hAC0;
        12'hE2E: sinewave <= 12'hAC3;
        12'hE2F: sinewave <= 12'hAC5;
        12'hE30: sinewave <= 12'hAC7;
        12'hE31: sinewave <= 12'hACA;
        12'hE32: sinewave <= 12'hACC;
        12'hE33: sinewave <= 12'hACF;
        12'hE34: sinewave <= 12'hAD1;
        12'hE35: sinewave <= 12'hAD3;
        12'hE36: sinewave <= 12'hAD6;
        12'hE37: sinewave <= 12'hAD8;
        12'hE38: sinewave <= 12'hADB;
        12'hE39: sinewave <= 12'hADD;
        12'hE3A: sinewave <= 12'hADF;
        12'hE3B: sinewave <= 12'hAE2;
        12'hE3C: sinewave <= 12'hAE4;
        12'hE3D: sinewave <= 12'hAE7;
        12'hE3E: sinewave <= 12'hAE9;
        12'hE3F: sinewave <= 12'hAEB;
        12'hE40: sinewave <= 12'hAEE;
        12'hE41: sinewave <= 12'hAF0;
        12'hE42: sinewave <= 12'hAF3;
        12'hE43: sinewave <= 12'hAF5;
        12'hE44: sinewave <= 12'hAF8;
        12'hE45: sinewave <= 12'hAFA;
        12'hE46: sinewave <= 12'hAFD;
        12'hE47: sinewave <= 12'hAFF;
        12'hE48: sinewave <= 12'hB01;
        12'hE49: sinewave <= 12'hB04;
        12'hE4A: sinewave <= 12'hB06;
        12'hE4B: sinewave <= 12'hB09;
        12'hE4C: sinewave <= 12'hB0B;
        12'hE4D: sinewave <= 12'hB0E;
        12'hE4E: sinewave <= 12'hB10;
        12'hE4F: sinewave <= 12'hB13;
        12'hE50: sinewave <= 12'hB15;
        12'hE51: sinewave <= 12'hB18;
        12'hE52: sinewave <= 12'hB1A;
        12'hE53: sinewave <= 12'hB1D;
        12'hE54: sinewave <= 12'hB1F;
        12'hE55: sinewave <= 12'hB22;
        12'hE56: sinewave <= 12'hB24;
        12'hE57: sinewave <= 12'hB27;
        12'hE58: sinewave <= 12'hB29;
        12'hE59: sinewave <= 12'hB2C;
        12'hE5A: sinewave <= 12'hB2E;
        12'hE5B: sinewave <= 12'hB31;
        12'hE5C: sinewave <= 12'hB33;
        12'hE5D: sinewave <= 12'hB36;
        12'hE5E: sinewave <= 12'hB38;
        12'hE5F: sinewave <= 12'hB3B;
        12'hE60: sinewave <= 12'hB3D;
        12'hE61: sinewave <= 12'hB40;
        12'hE62: sinewave <= 12'hB42;
        12'hE63: sinewave <= 12'hB45;
        12'hE64: sinewave <= 12'hB47;
        12'hE65: sinewave <= 12'hB4A;
        12'hE66: sinewave <= 12'hB4C;
        12'hE67: sinewave <= 12'hB4F;
        12'hE68: sinewave <= 12'hB51;
        12'hE69: sinewave <= 12'hB54;
        12'hE6A: sinewave <= 12'hB56;
        12'hE6B: sinewave <= 12'hB59;
        12'hE6C: sinewave <= 12'hB5C;
        12'hE6D: sinewave <= 12'hB5E;
        12'hE6E: sinewave <= 12'hB61;
        12'hE6F: sinewave <= 12'hB63;
        12'hE70: sinewave <= 12'hB66;
        12'hE71: sinewave <= 12'hB68;
        12'hE72: sinewave <= 12'hB6B;
        12'hE73: sinewave <= 12'hB6E;
        12'hE74: sinewave <= 12'hB70;
        12'hE75: sinewave <= 12'hB73;
        12'hE76: sinewave <= 12'hB75;
        12'hE77: sinewave <= 12'hB78;
        12'hE78: sinewave <= 12'hB7A;
        12'hE79: sinewave <= 12'hB7D;
        12'hE7A: sinewave <= 12'hB80;
        12'hE7B: sinewave <= 12'hB82;
        12'hE7C: sinewave <= 12'hB85;
        12'hE7D: sinewave <= 12'hB87;
        12'hE7E: sinewave <= 12'hB8A;
        12'hE7F: sinewave <= 12'hB8D;
        12'hE80: sinewave <= 12'hB8F;
        12'hE81: sinewave <= 12'hB92;
        12'hE82: sinewave <= 12'hB94;
        12'hE83: sinewave <= 12'hB97;
        12'hE84: sinewave <= 12'hB9A;
        12'hE85: sinewave <= 12'hB9C;
        12'hE86: sinewave <= 12'hB9F;
        12'hE87: sinewave <= 12'hBA2;
        12'hE88: sinewave <= 12'hBA4;
        12'hE89: sinewave <= 12'hBA7;
        12'hE8A: sinewave <= 12'hBA9;
        12'hE8B: sinewave <= 12'hBAC;
        12'hE8C: sinewave <= 12'hBAF;
        12'hE8D: sinewave <= 12'hBB1;
        12'hE8E: sinewave <= 12'hBB4;
        12'hE8F: sinewave <= 12'hBB7;
        12'hE90: sinewave <= 12'hBB9;
        12'hE91: sinewave <= 12'hBBC;
        12'hE92: sinewave <= 12'hBBF;
        12'hE93: sinewave <= 12'hBC1;
        12'hE94: sinewave <= 12'hBC4;
        12'hE95: sinewave <= 12'hBC7;
        12'hE96: sinewave <= 12'hBC9;
        12'hE97: sinewave <= 12'hBCC;
        12'hE98: sinewave <= 12'hBCF;
        12'hE99: sinewave <= 12'hBD1;
        12'hE9A: sinewave <= 12'hBD4;
        12'hE9B: sinewave <= 12'hBD7;
        12'hE9C: sinewave <= 12'hBD9;
        12'hE9D: sinewave <= 12'hBDC;
        12'hE9E: sinewave <= 12'hBDF;
        12'hE9F: sinewave <= 12'hBE1;
        12'hEA0: sinewave <= 12'hBE4;
        12'hEA1: sinewave <= 12'hBE7;
        12'hEA2: sinewave <= 12'hBEA;
        12'hEA3: sinewave <= 12'hBEC;
        12'hEA4: sinewave <= 12'hBEF;
        12'hEA5: sinewave <= 12'hBF2;
        12'hEA6: sinewave <= 12'hBF4;
        12'hEA7: sinewave <= 12'hBF7;
        12'hEA8: sinewave <= 12'hBFA;
        12'hEA9: sinewave <= 12'hBFC;
        12'hEAA: sinewave <= 12'hBFF;
        12'hEAB: sinewave <= 12'hC02;
        12'hEAC: sinewave <= 12'hC05;
        12'hEAD: sinewave <= 12'hC07;
        12'hEAE: sinewave <= 12'hC0A;
        12'hEAF: sinewave <= 12'hC0D;
        12'hEB0: sinewave <= 12'hC10;
        12'hEB1: sinewave <= 12'hC12;
        12'hEB2: sinewave <= 12'hC15;
        12'hEB3: sinewave <= 12'hC18;
        12'hEB4: sinewave <= 12'hC1A;
        12'hEB5: sinewave <= 12'hC1D;
        12'hEB6: sinewave <= 12'hC20;
        12'hEB7: sinewave <= 12'hC23;
        12'hEB8: sinewave <= 12'hC25;
        12'hEB9: sinewave <= 12'hC28;
        12'hEBA: sinewave <= 12'hC2B;
        12'hEBB: sinewave <= 12'hC2E;
        12'hEBC: sinewave <= 12'hC30;
        12'hEBD: sinewave <= 12'hC33;
        12'hEBE: sinewave <= 12'hC36;
        12'hEBF: sinewave <= 12'hC39;
        12'hEC0: sinewave <= 12'hC3C;
        12'hEC1: sinewave <= 12'hC3E;
        12'hEC2: sinewave <= 12'hC41;
        12'hEC3: sinewave <= 12'hC44;
        12'hEC4: sinewave <= 12'hC47;
        12'hEC5: sinewave <= 12'hC49;
        12'hEC6: sinewave <= 12'hC4C;
        12'hEC7: sinewave <= 12'hC4F;
        12'hEC8: sinewave <= 12'hC52;
        12'hEC9: sinewave <= 12'hC55;
        12'hECA: sinewave <= 12'hC57;
        12'hECB: sinewave <= 12'hC5A;
        12'hECC: sinewave <= 12'hC5D;
        12'hECD: sinewave <= 12'hC60;
        12'hECE: sinewave <= 12'hC63;
        12'hECF: sinewave <= 12'hC65;
        12'hED0: sinewave <= 12'hC68;
        12'hED1: sinewave <= 12'hC6B;
        12'hED2: sinewave <= 12'hC6E;
        12'hED3: sinewave <= 12'hC71;
        12'hED4: sinewave <= 12'hC73;
        12'hED5: sinewave <= 12'hC76;
        12'hED6: sinewave <= 12'hC79;
        12'hED7: sinewave <= 12'hC7C;
        12'hED8: sinewave <= 12'hC7F;
        12'hED9: sinewave <= 12'hC81;
        12'hEDA: sinewave <= 12'hC84;
        12'hEDB: sinewave <= 12'hC87;
        12'hEDC: sinewave <= 12'hC8A;
        12'hEDD: sinewave <= 12'hC8D;
        12'hEDE: sinewave <= 12'hC90;
        12'hEDF: sinewave <= 12'hC92;
        12'hEE0: sinewave <= 12'hC95;
        12'hEE1: sinewave <= 12'hC98;
        12'hEE2: sinewave <= 12'hC9B;
        12'hEE3: sinewave <= 12'hC9E;
        12'hEE4: sinewave <= 12'hCA1;
        12'hEE5: sinewave <= 12'hCA4;
        12'hEE6: sinewave <= 12'hCA6;
        12'hEE7: sinewave <= 12'hCA9;
        12'hEE8: sinewave <= 12'hCAC;
        12'hEE9: sinewave <= 12'hCAF;
        12'hEEA: sinewave <= 12'hCB2;
        12'hEEB: sinewave <= 12'hCB5;
        12'hEEC: sinewave <= 12'hCB8;
        12'hEED: sinewave <= 12'hCBA;
        12'hEEE: sinewave <= 12'hCBD;
        12'hEEF: sinewave <= 12'hCC0;
        12'hEF0: sinewave <= 12'hCC3;
        12'hEF1: sinewave <= 12'hCC6;
        12'hEF2: sinewave <= 12'hCC9;
        12'hEF3: sinewave <= 12'hCCC;
        12'hEF4: sinewave <= 12'hCCE;
        12'hEF5: sinewave <= 12'hCD1;
        12'hEF6: sinewave <= 12'hCD4;
        12'hEF7: sinewave <= 12'hCD7;
        12'hEF8: sinewave <= 12'hCDA;
        12'hEF9: sinewave <= 12'hCDD;
        12'hEFA: sinewave <= 12'hCE0;
        12'hEFB: sinewave <= 12'hCE3;
        12'hEFC: sinewave <= 12'hCE6;
        12'hEFD: sinewave <= 12'hCE8;
        12'hEFE: sinewave <= 12'hCEB;
        12'hEFF: sinewave <= 12'hCEE;
        12'hF00: sinewave <= 12'hCF1;
        12'hF01: sinewave <= 12'hCF4;
        12'hF02: sinewave <= 12'hCF7;
        12'hF03: sinewave <= 12'hCFA;
        12'hF04: sinewave <= 12'hCFD;
        12'hF05: sinewave <= 12'hD00;
        12'hF06: sinewave <= 12'hD03;
        12'hF07: sinewave <= 12'hD05;
        12'hF08: sinewave <= 12'hD08;
        12'hF09: sinewave <= 12'hD0B;
        12'hF0A: sinewave <= 12'hD0E;
        12'hF0B: sinewave <= 12'hD11;
        12'hF0C: sinewave <= 12'hD14;
        12'hF0D: sinewave <= 12'hD17;
        12'hF0E: sinewave <= 12'hD1A;
        12'hF0F: sinewave <= 12'hD1D;
        12'hF10: sinewave <= 12'hD20;
        12'hF11: sinewave <= 12'hD23;
        12'hF12: sinewave <= 12'hD26;
        12'hF13: sinewave <= 12'hD29;
        12'hF14: sinewave <= 12'hD2C;
        12'hF15: sinewave <= 12'hD2E;
        12'hF16: sinewave <= 12'hD31;
        12'hF17: sinewave <= 12'hD34;
        12'hF18: sinewave <= 12'hD37;
        12'hF19: sinewave <= 12'hD3A;
        12'hF1A: sinewave <= 12'hD3D;
        12'hF1B: sinewave <= 12'hD40;
        12'hF1C: sinewave <= 12'hD43;
        12'hF1D: sinewave <= 12'hD46;
        12'hF1E: sinewave <= 12'hD49;
        12'hF1F: sinewave <= 12'hD4C;
        12'hF20: sinewave <= 12'hD4F;
        12'hF21: sinewave <= 12'hD52;
        12'hF22: sinewave <= 12'hD55;
        12'hF23: sinewave <= 12'hD58;
        12'hF24: sinewave <= 12'hD5B;
        12'hF25: sinewave <= 12'hD5E;
        12'hF26: sinewave <= 12'hD61;
        12'hF27: sinewave <= 12'hD64;
        12'hF28: sinewave <= 12'hD67;
        12'hF29: sinewave <= 12'hD6A;
        12'hF2A: sinewave <= 12'hD6D;
        12'hF2B: sinewave <= 12'hD70;
        12'hF2C: sinewave <= 12'hD72;
        12'hF2D: sinewave <= 12'hD75;
        12'hF2E: sinewave <= 12'hD78;
        12'hF2F: sinewave <= 12'hD7B;
        12'hF30: sinewave <= 12'hD7E;
        12'hF31: sinewave <= 12'hD81;
        12'hF32: sinewave <= 12'hD84;
        12'hF33: sinewave <= 12'hD87;
        12'hF34: sinewave <= 12'hD8A;
        12'hF35: sinewave <= 12'hD8D;
        12'hF36: sinewave <= 12'hD90;
        12'hF37: sinewave <= 12'hD93;
        12'hF38: sinewave <= 12'hD96;
        12'hF39: sinewave <= 12'hD99;
        12'hF3A: sinewave <= 12'hD9C;
        12'hF3B: sinewave <= 12'hD9F;
        12'hF3C: sinewave <= 12'hDA2;
        12'hF3D: sinewave <= 12'hDA5;
        12'hF3E: sinewave <= 12'hDA8;
        12'hF3F: sinewave <= 12'hDAB;
        12'hF40: sinewave <= 12'hDAE;
        12'hF41: sinewave <= 12'hDB1;
        12'hF42: sinewave <= 12'hDB4;
        12'hF43: sinewave <= 12'hDB7;
        12'hF44: sinewave <= 12'hDBA;
        12'hF45: sinewave <= 12'hDBD;
        12'hF46: sinewave <= 12'hDC0;
        12'hF47: sinewave <= 12'hDC3;
        12'hF48: sinewave <= 12'hDC6;
        12'hF49: sinewave <= 12'hDC9;
        12'hF4A: sinewave <= 12'hDCC;
        12'hF4B: sinewave <= 12'hDCF;
        12'hF4C: sinewave <= 12'hDD2;
        12'hF4D: sinewave <= 12'hDD5;
        12'hF4E: sinewave <= 12'hDD8;
        12'hF4F: sinewave <= 12'hDDC;
        12'hF50: sinewave <= 12'hDDF;
        12'hF51: sinewave <= 12'hDE2;
        12'hF52: sinewave <= 12'hDE5;
        12'hF53: sinewave <= 12'hDE8;
        12'hF54: sinewave <= 12'hDEB;
        12'hF55: sinewave <= 12'hDEE;
        12'hF56: sinewave <= 12'hDF1;
        12'hF57: sinewave <= 12'hDF4;
        12'hF58: sinewave <= 12'hDF7;
        12'hF59: sinewave <= 12'hDFA;
        12'hF5A: sinewave <= 12'hDFD;
        12'hF5B: sinewave <= 12'hE00;
        12'hF5C: sinewave <= 12'hE03;
        12'hF5D: sinewave <= 12'hE06;
        12'hF5E: sinewave <= 12'hE09;
        12'hF5F: sinewave <= 12'hE0C;
        12'hF60: sinewave <= 12'hE0F;
        12'hF61: sinewave <= 12'hE12;
        12'hF62: sinewave <= 12'hE15;
        12'hF63: sinewave <= 12'hE18;
        12'hF64: sinewave <= 12'hE1B;
        12'hF65: sinewave <= 12'hE1E;
        12'hF66: sinewave <= 12'hE21;
        12'hF67: sinewave <= 12'hE24;
        12'hF68: sinewave <= 12'hE28;
        12'hF69: sinewave <= 12'hE2B;
        12'hF6A: sinewave <= 12'hE2E;
        12'hF6B: sinewave <= 12'hE31;
        12'hF6C: sinewave <= 12'hE34;
        12'hF6D: sinewave <= 12'hE37;
        12'hF6E: sinewave <= 12'hE3A;
        12'hF6F: sinewave <= 12'hE3D;
        12'hF70: sinewave <= 12'hE40;
        12'hF71: sinewave <= 12'hE43;
        12'hF72: sinewave <= 12'hE46;
        12'hF73: sinewave <= 12'hE49;
        12'hF74: sinewave <= 12'hE4C;
        12'hF75: sinewave <= 12'hE4F;
        12'hF76: sinewave <= 12'hE52;
        12'hF77: sinewave <= 12'hE55;
        12'hF78: sinewave <= 12'hE59;
        12'hF79: sinewave <= 12'hE5C;
        12'hF7A: sinewave <= 12'hE5F;
        12'hF7B: sinewave <= 12'hE62;
        12'hF7C: sinewave <= 12'hE65;
        12'hF7D: sinewave <= 12'hE68;
        12'hF7E: sinewave <= 12'hE6B;
        12'hF7F: sinewave <= 12'hE6E;
        12'hF80: sinewave <= 12'hE71;
        12'hF81: sinewave <= 12'hE74;
        12'hF82: sinewave <= 12'hE77;
        12'hF83: sinewave <= 12'hE7A;
        12'hF84: sinewave <= 12'hE7D;
        12'hF85: sinewave <= 12'hE81;
        12'hF86: sinewave <= 12'hE84;
        12'hF87: sinewave <= 12'hE87;
        12'hF88: sinewave <= 12'hE8A;
        12'hF89: sinewave <= 12'hE8D;
        12'hF8A: sinewave <= 12'hE90;
        12'hF8B: sinewave <= 12'hE93;
        12'hF8C: sinewave <= 12'hE96;
        12'hF8D: sinewave <= 12'hE99;
        12'hF8E: sinewave <= 12'hE9C;
        12'hF8F: sinewave <= 12'hE9F;
        12'hF90: sinewave <= 12'hEA3;
        12'hF91: sinewave <= 12'hEA6;
        12'hF92: sinewave <= 12'hEA9;
        12'hF93: sinewave <= 12'hEAC;
        12'hF94: sinewave <= 12'hEAF;
        12'hF95: sinewave <= 12'hEB2;
        12'hF96: sinewave <= 12'hEB5;
        12'hF97: sinewave <= 12'hEB8;
        12'hF98: sinewave <= 12'hEBB;
        12'hF99: sinewave <= 12'hEBE;
        12'hF9A: sinewave <= 12'hEC2;
        12'hF9B: sinewave <= 12'hEC5;
        12'hF9C: sinewave <= 12'hEC8;
        12'hF9D: sinewave <= 12'hECB;
        12'hF9E: sinewave <= 12'hECE;
        12'hF9F: sinewave <= 12'hED1;
        12'hFA0: sinewave <= 12'hED4;
        12'hFA1: sinewave <= 12'hED7;
        12'hFA2: sinewave <= 12'hEDA;
        12'hFA3: sinewave <= 12'hEDD;
        12'hFA4: sinewave <= 12'hEE1;
        12'hFA5: sinewave <= 12'hEE4;
        12'hFA6: sinewave <= 12'hEE7;
        12'hFA7: sinewave <= 12'hEEA;
        12'hFA8: sinewave <= 12'hEED;
        12'hFA9: sinewave <= 12'hEF0;
        12'hFAA: sinewave <= 12'hEF3;
        12'hFAB: sinewave <= 12'hEF6;
        12'hFAC: sinewave <= 12'hEF9;
        12'hFAD: sinewave <= 12'hEFD;
        12'hFAE: sinewave <= 12'hF00;
        12'hFAF: sinewave <= 12'hF03;
        12'hFB0: sinewave <= 12'hF06;
        12'hFB1: sinewave <= 12'hF09;
        12'hFB2: sinewave <= 12'hF0C;
        12'hFB3: sinewave <= 12'hF0F;
        12'hFB4: sinewave <= 12'hF12;
        12'hFB5: sinewave <= 12'hF16;
        12'hFB6: sinewave <= 12'hF19;
        12'hFB7: sinewave <= 12'hF1C;
        12'hFB8: sinewave <= 12'hF1F;
        12'hFB9: sinewave <= 12'hF22;
        12'hFBA: sinewave <= 12'hF25;
        12'hFBB: sinewave <= 12'hF28;
        12'hFBC: sinewave <= 12'hF2B;
        12'hFBD: sinewave <= 12'hF2E;
        12'hFBE: sinewave <= 12'hF32;
        12'hFBF: sinewave <= 12'hF35;
        12'hFC0: sinewave <= 12'hF38;
        12'hFC1: sinewave <= 12'hF3B;
        12'hFC2: sinewave <= 12'hF3E;
        12'hFC3: sinewave <= 12'hF41;
        12'hFC4: sinewave <= 12'hF44;
        12'hFC5: sinewave <= 12'hF47;
        12'hFC6: sinewave <= 12'hF4B;
        12'hFC7: sinewave <= 12'hF4E;
        12'hFC8: sinewave <= 12'hF51;
        12'hFC9: sinewave <= 12'hF54;
        12'hFCA: sinewave <= 12'hF57;
        12'hFCB: sinewave <= 12'hF5A;
        12'hFCC: sinewave <= 12'hF5D;
        12'hFCD: sinewave <= 12'hF61;
        12'hFCE: sinewave <= 12'hF64;
        12'hFCF: sinewave <= 12'hF67;
        12'hFD0: sinewave <= 12'hF6A;
        12'hFD1: sinewave <= 12'hF6D;
        12'hFD2: sinewave <= 12'hF70;
        12'hFD3: sinewave <= 12'hF73;
        12'hFD4: sinewave <= 12'hF76;
        12'hFD5: sinewave <= 12'hF7A;
        12'hFD6: sinewave <= 12'hF7D;
        12'hFD7: sinewave <= 12'hF80;
        12'hFD8: sinewave <= 12'hF83;
        12'hFD9: sinewave <= 12'hF86;
        12'hFDA: sinewave <= 12'hF89;
        12'hFDB: sinewave <= 12'hF8C;
        12'hFDC: sinewave <= 12'hF90;
        12'hFDD: sinewave <= 12'hF93;
        12'hFDE: sinewave <= 12'hF96;
        12'hFDF: sinewave <= 12'hF99;
        12'hFE0: sinewave <= 12'hF9C;
        12'hFE1: sinewave <= 12'hF9F;
        12'hFE2: sinewave <= 12'hFA2;
        12'hFE3: sinewave <= 12'hFA5;
        12'hFE4: sinewave <= 12'hFA9;
        12'hFE5: sinewave <= 12'hFAC;
        12'hFE6: sinewave <= 12'hFAF;
        12'hFE7: sinewave <= 12'hFB2;
        12'hFE8: sinewave <= 12'hFB5;
        12'hFE9: sinewave <= 12'hFB8;
        12'hFEA: sinewave <= 12'hFBB;
        12'hFEB: sinewave <= 12'hFBF;
        12'hFEC: sinewave <= 12'hFC2;
        12'hFED: sinewave <= 12'hFC5;
        12'hFEE: sinewave <= 12'hFC8;
        12'hFEF: sinewave <= 12'hFCB;
        12'hFF0: sinewave <= 12'hFCE;
        12'hFF1: sinewave <= 12'hFD1;
        12'hFF2: sinewave <= 12'hFD5;
        12'hFF3: sinewave <= 12'hFD8;
        12'hFF4: sinewave <= 12'hFDB;
        12'hFF5: sinewave <= 12'hFDE;
        12'hFF6: sinewave <= 12'hFE1;
        12'hFF7: sinewave <= 12'hFE4;
        12'hFF8: sinewave <= 12'hFE7;
        12'hFF9: sinewave <= 12'hFEB;
        12'hFFA: sinewave <= 12'hFEE;
        12'hFFB: sinewave <= 12'hFF1;
        12'hFFC: sinewave <= 12'hFF4;
        12'hFFD: sinewave <= 12'hFF7;
        12'hFFE: sinewave <= 12'hFFA;
        12'hFFF: sinewave <= 12'hFFD;
        endcase
    end
end

initial begin
	$dumpfile("simpleSine_waves.vcd");
	$dumpvars;
end

endmodule